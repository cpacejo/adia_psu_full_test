magic
tech sky130A
magscale 1 2
timestamp 1717221846
<< metal3 >>
rect -9798 2812 -3426 2840
rect -9798 -2812 -3510 2812
rect -3446 -2812 -3426 2812
rect -9798 -2840 -3426 -2812
rect -3186 2812 3186 2840
rect -3186 -2812 3102 2812
rect 3166 -2812 3186 2812
rect -3186 -2840 3186 -2812
rect 3426 2812 9798 2840
rect 3426 -2812 9714 2812
rect 9778 -2812 9798 2812
rect 3426 -2840 9798 -2812
<< via3 >>
rect -3510 -2812 -3446 2812
rect 3102 -2812 3166 2812
rect 9714 -2812 9778 2812
<< mimcap >>
rect -9758 2760 -3758 2800
rect -9758 -2760 -9718 2760
rect -3798 -2760 -3758 2760
rect -9758 -2800 -3758 -2760
rect -3146 2760 2854 2800
rect -3146 -2760 -3106 2760
rect 2814 -2760 2854 2760
rect -3146 -2800 2854 -2760
rect 3466 2760 9466 2800
rect 3466 -2760 3506 2760
rect 9426 -2760 9466 2760
rect 3466 -2800 9466 -2760
<< mimcapcontact >>
rect -9718 -2760 -3798 2760
rect -3106 -2760 2814 2760
rect 3506 -2760 9426 2760
<< metal4 >>
rect -3526 2812 -3430 2828
rect -9719 2760 -3797 2761
rect -9719 -2760 -9718 2760
rect -3798 -2760 -3797 2760
rect -9719 -2761 -3797 -2760
rect -3526 -2812 -3510 2812
rect -3446 -2812 -3430 2812
rect 3086 2812 3182 2828
rect -3107 2760 2815 2761
rect -3107 -2760 -3106 2760
rect 2814 -2760 2815 2760
rect -3107 -2761 2815 -2760
rect -3526 -2828 -3430 -2812
rect 3086 -2812 3102 2812
rect 3166 -2812 3182 2812
rect 9698 2812 9794 2828
rect 3505 2760 9427 2761
rect 3505 -2760 3506 2760
rect 9426 -2760 9427 2760
rect 3505 -2761 9427 -2760
rect 3086 -2828 3182 -2812
rect 9698 -2812 9714 2812
rect 9778 -2812 9794 2812
rect 9698 -2828 9794 -2812
<< properties >>
string FIXED_BBOX 3426 -2840 9506 2840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 28 val 1.702k carea 2.00 cperi 0.19 nx 3 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
