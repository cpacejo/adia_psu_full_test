magic
tech sky130A
magscale 1 2
timestamp 1717221846
<< error_s >>
rect 4086 22370 4144 22376
rect 4086 22336 4098 22370
rect 4086 22330 4144 22336
rect 4086 22176 4144 22182
rect 3174 22158 3232 22164
rect 3174 22124 3186 22158
rect 4086 22142 4098 22176
rect 4086 22136 4144 22142
rect 3174 22118 3232 22124
rect 3174 21830 3232 21836
rect 3174 21796 3186 21830
rect 3174 21790 3232 21796
<< locali >>
rect 11640 37580 11920 37660
rect 11660 37020 11880 37080
rect 11640 31580 11920 31660
rect 11660 31020 11880 31080
rect 11640 25580 11920 25660
rect 11660 25020 11880 25080
rect 11640 19580 11920 19660
rect 11660 19020 11880 19080
rect 11640 13580 11920 13660
rect 11660 13020 11880 13080
rect 11640 7580 11920 7660
rect 11660 7020 11880 7080
rect 11640 1580 11920 1660
rect 11660 1020 11880 1080
<< viali >>
rect 11470 37336 11506 37371
rect 11562 37317 11608 37363
rect 11470 31336 11506 31371
rect 11562 31317 11608 31363
rect 11468 25336 11504 25371
rect 11562 25317 11608 25363
rect 11468 19335 11507 19374
rect 11562 19337 11608 19383
rect 11469 13336 11505 13371
rect 11562 13317 11608 13363
rect 11470 7337 11506 7372
rect 11562 7317 11608 7363
rect 11468 1336 11504 1371
rect 11562 1317 11608 1363
<< metal1 >>
rect 11670 44490 11730 44496
rect 11210 44430 11670 44490
rect 9590 43890 9650 43896
rect 10270 43890 10330 43896
rect 9650 43830 10270 43890
rect 9590 43824 9650 43830
rect 10270 43824 10330 43830
rect 11210 42850 11270 44430
rect 11670 44424 11730 44430
rect 11210 42784 11270 42790
rect 11050 42630 11110 42636
rect 9424 42570 9430 42630
rect 9490 42570 11050 42630
rect 11050 42564 11110 42570
rect 10850 42410 10910 42416
rect 9424 42350 9430 42410
rect 9490 42350 10850 42410
rect 10850 42344 10910 42350
rect 10650 39010 10710 39016
rect 9504 38950 9510 39010
rect 9570 38950 10650 39010
rect 10650 38944 10710 38950
rect 11773 38101 11779 38161
rect 11839 38101 11845 38161
rect 11779 37820 11839 38101
rect 11240 37760 12160 37820
rect 11240 37380 11300 37760
rect 12080 37740 12160 37760
rect 11998 37710 12044 37722
rect 11998 37704 12004 37710
rect 11996 37676 12036 37704
rect 12038 37676 12044 37710
rect 11996 37664 12044 37676
rect 12192 37710 12238 37722
rect 12192 37704 12198 37710
rect 12232 37704 12238 37710
rect 12192 37664 12238 37704
rect 11800 37540 11900 37560
rect 11800 37480 11820 37540
rect 11880 37494 11900 37540
rect 11996 37494 12036 37664
rect 11880 37480 12036 37494
rect 11800 37460 12036 37480
rect 11836 37454 12036 37460
rect 12196 37494 12236 37664
rect 12360 37520 12460 37540
rect 12360 37494 12380 37520
rect 12196 37460 12380 37494
rect 12440 37460 12460 37520
rect 12196 37454 12460 37460
rect 11240 37371 11520 37380
rect 11240 37340 11470 37371
rect 11250 37336 11470 37340
rect 11506 37336 11520 37371
rect 11250 37330 11520 37336
rect 11556 37363 11614 37375
rect 11556 37317 11562 37363
rect 11608 37317 11763 37363
rect 11556 37305 11614 37317
rect 11717 37163 11763 37317
rect 11836 37262 11876 37454
rect 12360 37440 12460 37454
rect 12366 37262 12406 37440
rect 11832 37214 11878 37262
rect 11832 37212 11838 37214
rect 11872 37212 11878 37214
rect 11832 37200 11878 37212
rect 12360 37214 12406 37262
rect 12360 37212 12366 37214
rect 12400 37212 12406 37214
rect 12360 37200 12406 37212
rect 11717 37117 11963 37163
rect 10470 34930 10530 34936
rect 9564 34870 9570 34930
rect 9630 34870 10470 34930
rect 10470 34864 10530 34870
rect 10090 33390 10150 33396
rect 8764 33330 8770 33390
rect 8830 33330 10090 33390
rect 10090 33324 10150 33330
rect 11200 32690 11280 32700
rect 9544 32630 9550 32690
rect 9610 32630 11210 32690
rect 11270 32630 11280 32690
rect 11200 32620 11280 32630
rect 11726 32027 11732 32087
rect 11792 32027 11798 32087
rect 11732 31820 11792 32027
rect 11240 31760 12160 31820
rect 11240 31380 11300 31760
rect 11732 31752 11792 31760
rect 12080 31740 12160 31760
rect 11998 31710 12044 31722
rect 11998 31704 12004 31710
rect 11996 31676 12036 31704
rect 12038 31676 12044 31710
rect 11996 31664 12044 31676
rect 12192 31710 12238 31722
rect 12192 31704 12198 31710
rect 12232 31704 12238 31710
rect 12192 31664 12238 31704
rect 11800 31540 11900 31560
rect 11800 31480 11820 31540
rect 11880 31494 11900 31540
rect 11996 31494 12036 31664
rect 11880 31480 12036 31494
rect 11800 31460 12036 31480
rect 11836 31454 12036 31460
rect 12196 31494 12236 31664
rect 12360 31520 12460 31540
rect 12360 31494 12380 31520
rect 12196 31460 12380 31494
rect 12440 31460 12460 31520
rect 12196 31454 12460 31460
rect 11240 31371 11520 31380
rect 11240 31340 11470 31371
rect 11250 31336 11470 31340
rect 11506 31336 11520 31371
rect 11250 31330 11520 31336
rect 11556 31363 11614 31375
rect 11556 31317 11562 31363
rect 11608 31317 11763 31363
rect 11556 31305 11614 31317
rect 11717 31163 11763 31317
rect 11836 31262 11876 31454
rect 12360 31440 12460 31454
rect 12366 31262 12406 31440
rect 11832 31214 11878 31262
rect 11832 31212 11838 31214
rect 11872 31212 11878 31214
rect 11832 31200 11878 31212
rect 12360 31214 12406 31262
rect 12360 31212 12366 31214
rect 12400 31212 12406 31214
rect 12360 31200 12406 31212
rect 11717 31117 11983 31163
rect 11240 25810 12160 25820
rect 11240 25760 11688 25810
rect 11240 25380 11300 25760
rect 11598 25750 11688 25760
rect 11748 25760 12160 25810
rect 11748 25750 11754 25760
rect 12080 25740 12160 25760
rect 11998 25710 12044 25722
rect 11998 25704 12004 25710
rect 11996 25676 12036 25704
rect 12038 25676 12044 25710
rect 11996 25664 12044 25676
rect 12192 25710 12238 25722
rect 12192 25704 12198 25710
rect 12232 25704 12238 25710
rect 12192 25664 12238 25704
rect 11800 25540 11900 25560
rect 11800 25480 11820 25540
rect 11880 25494 11900 25540
rect 11996 25494 12036 25664
rect 11880 25480 12036 25494
rect 11800 25460 12036 25480
rect 11836 25454 12036 25460
rect 12196 25494 12236 25664
rect 12360 25520 12460 25540
rect 12360 25494 12380 25520
rect 12196 25460 12380 25494
rect 12440 25460 12460 25520
rect 12196 25454 12460 25460
rect 11240 25371 11520 25380
rect 11240 25340 11468 25371
rect 11250 25336 11468 25340
rect 11504 25336 11520 25371
rect 11250 25330 11520 25336
rect 11556 25363 11614 25375
rect 11556 25317 11562 25363
rect 11608 25317 11743 25363
rect 11556 25305 11614 25317
rect 11697 25163 11743 25317
rect 11836 25262 11876 25454
rect 12360 25440 12460 25454
rect 12366 25262 12406 25440
rect 11832 25214 11878 25262
rect 11832 25212 11838 25214
rect 11872 25212 11878 25214
rect 11832 25200 11878 25212
rect 12360 25214 12406 25262
rect 12360 25212 12366 25214
rect 12400 25212 12406 25214
rect 12360 25200 12406 25212
rect 11697 25117 11983 25163
rect 2730 23540 3010 23580
rect 2730 23410 2770 23540
rect 2520 23370 2770 23410
rect 2520 23170 2770 23210
rect 2730 23050 2770 23170
rect 2730 23010 3010 23050
rect 11559 19888 11565 19948
rect 11625 19888 11631 19948
rect 11565 19820 11625 19888
rect 11240 19760 12160 19820
rect 11240 19380 11300 19760
rect 12080 19740 12160 19760
rect 11998 19710 12044 19722
rect 11998 19704 12004 19710
rect 11996 19676 12036 19704
rect 12038 19676 12044 19710
rect 11996 19664 12044 19676
rect 12192 19710 12238 19722
rect 12192 19704 12198 19710
rect 12232 19704 12238 19710
rect 12192 19664 12238 19704
rect 11800 19540 11900 19560
rect 11800 19480 11820 19540
rect 11880 19494 11900 19540
rect 11996 19494 12036 19664
rect 11880 19480 12036 19494
rect 11800 19460 12036 19480
rect 11836 19454 12036 19460
rect 12196 19494 12236 19664
rect 12360 19520 12460 19540
rect 12360 19494 12380 19520
rect 12196 19460 12380 19494
rect 12440 19460 12460 19520
rect 12196 19454 12460 19460
rect 11556 19383 11614 19395
rect 11240 19374 11520 19380
rect 11240 19340 11468 19374
rect 11250 19335 11468 19340
rect 11507 19335 11520 19374
rect 11250 19330 11520 19335
rect 11556 19337 11562 19383
rect 11608 19337 11763 19383
rect 11460 19326 11515 19330
rect 11556 19325 11614 19337
rect 11717 19163 11763 19337
rect 11836 19262 11876 19454
rect 12360 19440 12460 19454
rect 12366 19262 12406 19440
rect 11832 19214 11878 19262
rect 11832 19212 11838 19214
rect 11872 19212 11878 19214
rect 11832 19200 11878 19212
rect 12360 19214 12406 19262
rect 12360 19212 12366 19214
rect 12400 19212 12406 19214
rect 12360 19200 12406 19212
rect 11717 19117 11963 19163
rect 11734 13858 11740 13918
rect 11800 13858 11806 13918
rect 11740 13820 11800 13858
rect 11240 13760 12160 13820
rect 11240 13380 11300 13760
rect 11740 13755 11800 13760
rect 12080 13740 12160 13760
rect 11998 13710 12044 13722
rect 11998 13704 12004 13710
rect 11996 13676 12036 13704
rect 12038 13676 12044 13710
rect 11996 13664 12044 13676
rect 12192 13710 12238 13722
rect 12192 13704 12198 13710
rect 12232 13704 12238 13710
rect 12192 13664 12238 13704
rect 11760 13540 11860 13560
rect 11760 13480 11780 13540
rect 11840 13494 11860 13540
rect 11996 13494 12036 13664
rect 11840 13480 12036 13494
rect 11760 13460 12036 13480
rect 11836 13454 12036 13460
rect 12196 13494 12236 13664
rect 12360 13520 12460 13540
rect 12360 13494 12380 13520
rect 12196 13460 12380 13494
rect 12440 13460 12460 13520
rect 12196 13454 12460 13460
rect 11240 13371 11520 13380
rect 11240 13340 11469 13371
rect 11250 13336 11469 13340
rect 11505 13336 11520 13371
rect 11250 13330 11520 13336
rect 11556 13363 11614 13375
rect 11556 13317 11562 13363
rect 11608 13317 11703 13363
rect 11556 13305 11614 13317
rect 11657 13183 11703 13317
rect 11836 13262 11876 13454
rect 12360 13440 12460 13454
rect 12366 13262 12406 13440
rect 11832 13214 11878 13262
rect 11832 13212 11838 13214
rect 11872 13212 11878 13214
rect 11832 13200 11878 13212
rect 12360 13214 12406 13262
rect 12360 13212 12366 13214
rect 12400 13212 12406 13214
rect 12360 13200 12406 13212
rect 11657 13143 11763 13183
rect 11917 13143 11963 13183
rect 11657 13137 11963 13143
rect 11717 13097 11963 13137
rect 11566 7908 11572 7968
rect 11632 7908 11638 7968
rect 11572 7820 11632 7908
rect 11240 7760 12160 7820
rect 11240 7380 11300 7760
rect 11998 7710 12044 7722
rect 12080 7720 12160 7760
rect 11998 7704 12004 7710
rect 11996 7676 12036 7704
rect 12038 7676 12044 7710
rect 11996 7664 12044 7676
rect 12192 7710 12238 7722
rect 12192 7704 12198 7710
rect 12232 7704 12238 7710
rect 12192 7664 12238 7704
rect 11760 7540 11860 7560
rect 11760 7480 11780 7540
rect 11840 7494 11860 7540
rect 11996 7494 12036 7664
rect 11840 7480 12036 7494
rect 11760 7460 12036 7480
rect 11836 7454 12036 7460
rect 12196 7494 12236 7664
rect 12360 7520 12460 7540
rect 12360 7494 12380 7520
rect 12196 7460 12380 7494
rect 12440 7460 12460 7520
rect 12196 7454 12460 7460
rect 11240 7372 11520 7380
rect 11240 7340 11470 7372
rect 11250 7337 11470 7340
rect 11506 7337 11520 7372
rect 11250 7330 11520 7337
rect 11556 7363 11614 7375
rect 11556 7317 11562 7363
rect 11608 7317 11703 7363
rect 11556 7305 11614 7317
rect 11657 7183 11703 7317
rect 11836 7262 11876 7454
rect 12360 7440 12460 7454
rect 12366 7262 12406 7440
rect 11832 7214 11878 7262
rect 11832 7212 11838 7214
rect 11872 7212 11878 7214
rect 11832 7200 11878 7212
rect 12360 7214 12406 7262
rect 12360 7212 12366 7214
rect 12400 7212 12406 7214
rect 12360 7200 12406 7212
rect 11657 7143 11783 7183
rect 11917 7143 11963 7183
rect 11657 7137 11963 7143
rect 11737 7097 11963 7137
rect 11369 1954 11375 2014
rect 11435 1954 11441 2014
rect 11375 1820 11435 1954
rect 11240 1760 12160 1820
rect 11240 1380 11300 1760
rect 11375 1752 11435 1760
rect 11998 1710 12044 1722
rect 11998 1704 12004 1710
rect 11996 1676 12036 1704
rect 12038 1676 12044 1710
rect 11996 1664 12044 1676
rect 12192 1710 12238 1722
rect 12192 1704 12198 1710
rect 12232 1704 12238 1710
rect 12192 1664 12238 1704
rect 11760 1540 11860 1560
rect 11760 1480 11780 1540
rect 11840 1494 11860 1540
rect 11996 1494 12036 1664
rect 11840 1480 12036 1494
rect 11760 1460 12036 1480
rect 11836 1454 12036 1460
rect 12196 1494 12236 1664
rect 12360 1520 12460 1540
rect 12360 1494 12380 1520
rect 12196 1460 12380 1494
rect 12440 1460 12460 1520
rect 12196 1454 12460 1460
rect 11240 1371 11520 1380
rect 11240 1340 11468 1371
rect 11250 1336 11468 1340
rect 11504 1336 11520 1371
rect 11250 1330 11520 1336
rect 11556 1363 11614 1375
rect 11556 1317 11562 1363
rect 11608 1358 11614 1363
rect 11608 1322 11698 1358
rect 11608 1317 11614 1322
rect 11556 1305 11614 1317
rect 11662 1178 11698 1322
rect 11836 1262 11876 1454
rect 12360 1440 12460 1454
rect 12366 1262 12406 1440
rect 11832 1214 11878 1262
rect 11832 1212 11838 1214
rect 11872 1212 11878 1214
rect 11832 1200 11878 1212
rect 12360 1214 12406 1262
rect 12360 1212 12366 1214
rect 12400 1212 12406 1214
rect 12360 1200 12406 1212
rect 11662 1158 11798 1178
rect 11662 1142 11978 1158
rect 11762 1122 11978 1142
<< via1 >>
rect 11670 44430 11730 44490
rect 9590 43830 9650 43890
rect 10270 43830 10330 43890
rect 11210 42790 11270 42850
rect 9430 42570 9490 42630
rect 11050 42570 11110 42630
rect 9430 42350 9490 42410
rect 10850 42350 10910 42410
rect 9510 38950 9570 39010
rect 10650 38950 10710 39010
rect 11779 38101 11839 38161
rect 11820 37480 11880 37540
rect 12380 37460 12440 37520
rect 9570 34870 9630 34930
rect 10470 34870 10530 34930
rect 8770 33330 8830 33390
rect 10090 33330 10150 33390
rect 9550 32630 9610 32690
rect 11210 32630 11270 32690
rect 11732 32027 11792 32087
rect 11820 31480 11880 31540
rect 12380 31460 12440 31520
rect 11688 25750 11748 25810
rect 11820 25480 11880 25540
rect 12380 25460 12440 25520
rect 11565 19888 11625 19948
rect 11820 19480 11880 19540
rect 12380 19460 12440 19520
rect 11740 13858 11800 13918
rect 11780 13480 11840 13540
rect 12380 13460 12440 13520
rect 11572 7908 11632 7968
rect 11780 7480 11840 7540
rect 12380 7460 12440 7520
rect 11375 1954 11435 2014
rect 11780 1480 11840 1540
rect 12380 1460 12440 1520
<< metal2 >>
rect 9350 44768 9410 44770
rect 9343 44712 9352 44768
rect 9408 44712 9417 44768
rect 6632 44150 6688 44157
rect 6370 44148 6690 44150
rect 6370 44092 6632 44148
rect 6688 44092 6690 44148
rect 6370 44090 6690 44092
rect 8294 44140 8354 44149
rect 6632 44083 6688 44090
rect 8294 44071 8354 44080
rect 3150 43728 3210 43910
rect 3143 43672 3152 43728
rect 3208 43672 3217 43728
rect 3150 43670 3210 43672
rect 9350 43650 9410 44712
rect 24350 44657 24410 44659
rect 12574 44628 12634 44630
rect 14046 44628 14106 44630
rect 14782 44628 14842 44630
rect 11838 44608 11898 44610
rect 9752 44590 9808 44597
rect 9750 44588 9810 44590
rect 9750 44532 9752 44588
rect 9808 44532 9810 44588
rect 11831 44552 11840 44608
rect 11896 44552 11905 44608
rect 12567 44572 12576 44628
rect 12632 44572 12641 44628
rect 13310 44608 13370 44610
rect 9584 43830 9590 43890
rect 9650 43830 9656 43890
rect 9590 43670 9650 43830
rect 9350 43581 9410 43590
rect 9430 42630 9490 42636
rect 9121 42570 9130 42630
rect 9190 42570 9430 42630
rect 9430 42564 9490 42570
rect 9430 42410 9490 42416
rect 9281 42350 9290 42410
rect 9350 42350 9430 42410
rect 9430 42344 9490 42350
rect 9510 39010 9570 39016
rect 9361 38950 9370 39010
rect 9430 38950 9510 39010
rect 9510 38944 9570 38950
rect 941 37610 950 37670
rect 1010 37610 1019 37670
rect 761 34210 770 34270
rect 830 34210 839 34270
rect 770 32310 830 34210
rect 950 32490 1010 37610
rect 1121 36230 1130 36290
rect 1190 36230 1199 36290
rect 1130 32690 1190 36230
rect 9570 34930 9630 34936
rect 9421 34870 9430 34930
rect 9490 34870 9570 34930
rect 9570 34864 9630 34870
rect 9350 33988 9410 33990
rect 9343 33932 9352 33988
rect 9408 33932 9417 33988
rect 8770 33390 8830 33396
rect 7010 33330 8770 33390
rect 8770 33324 8830 33330
rect 5472 33190 5528 33197
rect 9350 33190 9410 33932
rect 5470 33188 5770 33190
rect 5470 33132 5472 33188
rect 5528 33132 5770 33188
rect 5470 33130 5770 33132
rect 8950 33130 9410 33190
rect 5472 33123 5528 33130
rect 9550 32690 9610 32696
rect 1130 32630 9550 32690
rect 9550 32624 9610 32630
rect 9750 32490 9810 44532
rect 11838 44490 11898 44552
rect 11664 44430 11670 44490
rect 11730 44430 11898 44490
rect 12574 44330 12634 44572
rect 13303 44552 13312 44608
rect 13368 44552 13377 44608
rect 14039 44572 14048 44628
rect 14104 44572 14113 44628
rect 14775 44572 14784 44628
rect 14840 44572 14849 44628
rect 15518 44608 15578 44610
rect 16254 44608 16314 44610
rect 9950 44320 12634 44330
rect 9920 44270 12634 44320
rect 9920 32490 9980 44270
rect 13310 44110 13370 44552
rect 10090 44050 13370 44110
rect 10090 33390 10150 44050
rect 14046 43890 14106 44572
rect 10264 43830 10270 43890
rect 10330 43830 14106 43890
rect 10084 33330 10090 33390
rect 10150 33330 10156 33390
rect 950 32430 9980 32490
rect 9750 32310 9810 32430
rect 770 32250 9810 32310
rect 9750 32170 9810 32250
rect 9920 32200 9980 32430
rect 10090 32210 10150 33330
rect 10270 32210 10330 43830
rect 14782 43690 14842 44572
rect 15511 44552 15520 44608
rect 15576 44552 15585 44608
rect 16247 44552 16256 44608
rect 16312 44552 16321 44608
rect 24343 44601 24352 44657
rect 24408 44601 24417 44657
rect 16990 44568 17050 44570
rect 10470 43630 14842 43690
rect 10470 34930 10530 43630
rect 15518 43490 15578 44552
rect 10650 43430 15578 43490
rect 10650 39010 10710 43430
rect 16254 43290 16314 44552
rect 16983 44512 16992 44568
rect 17048 44512 17057 44568
rect 10850 43230 16314 43290
rect 10850 42410 10910 43230
rect 16990 43110 17050 44512
rect 11050 43050 17050 43110
rect 11050 42630 11110 43050
rect 24350 42862 24410 44601
rect 11204 42790 11210 42850
rect 11270 42790 11276 42850
rect 11375 42802 24410 42862
rect 11044 42570 11050 42630
rect 11110 42570 11116 42630
rect 10844 42350 10850 42410
rect 10910 42350 10916 42410
rect 10644 38950 10650 39010
rect 10710 38950 10716 39010
rect 10464 34870 10470 34930
rect 10530 34870 10536 34930
rect 10470 32230 10530 34870
rect 10650 32230 10710 38950
rect 10850 32230 10910 42350
rect 11050 32230 11110 42570
rect 11210 32690 11270 42790
rect 11375 42664 11435 42802
rect 11375 42595 11435 42604
rect 11779 38161 11839 38167
rect 12082 38161 12138 38168
rect 11839 38159 12140 38161
rect 11839 38103 12082 38159
rect 12138 38103 12140 38159
rect 11839 38101 12140 38103
rect 11779 38095 11839 38101
rect 12082 38094 12138 38101
rect 11800 37540 11900 37560
rect 11800 37480 11820 37540
rect 11880 37480 11900 37540
rect 11800 37286 11900 37480
rect 12360 37520 12460 37540
rect 12360 37460 12380 37520
rect 12440 37460 12460 37520
rect 12360 37440 12460 37460
rect 11800 37280 11902 37286
rect 11821 36923 11902 37280
rect 11821 36842 12149 36923
rect 11210 32230 11270 32630
rect 11732 32087 11792 32093
rect 11890 32087 11946 32094
rect 11792 32085 11948 32087
rect 11792 32029 11890 32085
rect 11946 32029 11948 32085
rect 11792 32027 11948 32029
rect 11732 32021 11792 32027
rect 11890 32020 11946 32027
rect 12068 31839 12149 36842
rect 11813 31758 12149 31839
rect 11813 31540 11894 31758
rect 11813 31480 11820 31540
rect 11880 31480 11894 31540
rect 11688 26055 11748 26057
rect 11681 25999 11690 26055
rect 11746 25999 11755 26055
rect 11688 25810 11748 25999
rect 11688 25744 11748 25750
rect 11813 25540 11894 31480
rect 12360 31520 12460 31540
rect 12360 31460 12380 31520
rect 12440 31460 12460 31520
rect 12360 31440 12460 31460
rect 11813 25480 11820 25540
rect 11880 25480 11894 25540
rect 11565 20099 11625 20101
rect 11558 20043 11567 20099
rect 11623 20043 11632 20099
rect 11565 19948 11625 20043
rect 11565 19882 11625 19888
rect 11813 19540 11894 25480
rect 12360 25520 12460 25540
rect 12360 25460 12380 25520
rect 12440 25460 12460 25520
rect 12360 25440 12460 25460
rect 11813 19480 11820 19540
rect 11880 19480 11894 19540
rect 11813 18939 11894 19480
rect 12360 19520 12460 19540
rect 12360 19460 12380 19520
rect 12440 19460 12460 19520
rect 12360 19440 12460 19460
rect 11813 18858 11953 18939
rect 11740 14049 11800 14051
rect 11733 13993 11742 14049
rect 11798 13993 11807 14049
rect 11740 13918 11800 13993
rect 11740 13852 11800 13858
rect 11872 13730 11953 18858
rect 11765 13649 11953 13730
rect 11765 13540 11846 13649
rect 11765 13480 11780 13540
rect 11840 13480 11846 13540
rect 11572 8130 11632 8132
rect 11565 8074 11574 8130
rect 11630 8074 11639 8130
rect 11572 7968 11632 8074
rect 11572 7902 11632 7908
rect 11765 7540 11846 13480
rect 12360 13520 12460 13540
rect 12360 13460 12380 13520
rect 12440 13460 12460 13520
rect 12360 13440 12460 13460
rect 11765 7480 11780 7540
rect 11840 7480 11846 7540
rect 11375 2233 11435 2235
rect 11368 2177 11377 2233
rect 11433 2177 11442 2233
rect 11375 2014 11435 2177
rect 11375 1948 11435 1954
rect 11765 1560 11846 7480
rect 12360 7520 12460 7540
rect 12360 7460 12380 7520
rect 12440 7460 12460 7520
rect 12360 7440 12460 7460
rect 11760 1540 11860 1560
rect 11760 1480 11780 1540
rect 11840 1480 11860 1540
rect 11760 830 11860 1480
rect 12360 1520 12460 1540
rect 12360 1460 12380 1520
rect 12440 1460 12460 1520
rect 12360 1440 12460 1460
rect 30515 830 30685 834
rect 11760 825 30690 830
rect 11760 800 30515 825
rect 11770 655 30515 800
rect 30685 655 30690 825
rect 11770 650 30690 655
rect 30515 646 30685 650
<< via2 >>
rect 9352 44712 9408 44768
rect 6632 44092 6688 44148
rect 8294 44080 8354 44140
rect 3152 43672 3208 43728
rect 9752 44532 9808 44588
rect 11840 44552 11896 44608
rect 12576 44572 12632 44628
rect 9350 43590 9410 43650
rect 9130 42570 9190 42630
rect 9290 42350 9350 42410
rect 9370 38950 9430 39010
rect 950 37610 1010 37670
rect 770 34210 830 34270
rect 1130 36230 1190 36290
rect 9430 34870 9490 34930
rect 9352 33932 9408 33988
rect 5472 33132 5528 33188
rect 13312 44552 13368 44608
rect 14048 44572 14104 44628
rect 14784 44572 14840 44628
rect 15520 44552 15576 44608
rect 16256 44552 16312 44608
rect 24352 44601 24408 44657
rect 16992 44512 17048 44568
rect 11375 42604 11435 42664
rect 12082 38103 12138 38159
rect 12380 37460 12440 37520
rect 11890 32029 11946 32085
rect 11690 25999 11746 26055
rect 12380 31460 12440 31520
rect 11567 20043 11623 20099
rect 12380 25460 12440 25520
rect 12380 19460 12440 19520
rect 11742 13993 11798 14049
rect 11574 8074 11630 8130
rect 12380 13460 12440 13520
rect 11377 2177 11433 2233
rect 12380 7460 12440 7520
rect 12380 1460 12440 1520
rect 30515 655 30685 825
<< metal3 >>
rect 9347 44770 9413 44773
rect 10364 44772 10428 44778
rect 9347 44768 10364 44770
rect 8156 44752 8220 44758
rect 390 44690 8156 44750
rect 390 33190 450 44690
rect 9347 44712 9352 44768
rect 9408 44712 10364 44768
rect 9347 44710 10364 44712
rect 9347 44707 9413 44710
rect 11094 44728 11100 44792
rect 11164 44728 11170 44792
rect 11830 44728 11836 44792
rect 11900 44728 11906 44792
rect 12566 44748 12572 44812
rect 12636 44748 12642 44812
rect 13302 44748 13308 44812
rect 13372 44748 13378 44812
rect 14038 44748 14044 44812
rect 14108 44748 14114 44812
rect 10364 44702 10428 44708
rect 8156 44682 8220 44688
rect 988 44592 1052 44598
rect 610 44530 988 44590
rect 610 43050 670 44530
rect 988 44522 1052 44528
rect 9747 44590 9813 44593
rect 11102 44590 11162 44728
rect 11838 44613 11898 44728
rect 12574 44633 12634 44748
rect 12571 44628 12637 44633
rect 9747 44588 11162 44590
rect 9747 44532 9752 44588
rect 9808 44532 11162 44588
rect 11835 44608 11901 44613
rect 11835 44552 11840 44608
rect 11896 44552 11901 44608
rect 12571 44572 12576 44628
rect 12632 44572 12637 44628
rect 13310 44613 13370 44748
rect 14046 44633 14106 44748
rect 14774 44728 14780 44792
rect 14844 44728 14850 44792
rect 15510 44748 15516 44812
rect 15580 44748 15586 44812
rect 14782 44633 14842 44728
rect 14043 44628 14109 44633
rect 12571 44567 12637 44572
rect 13307 44608 13373 44613
rect 11835 44547 11901 44552
rect 13307 44552 13312 44608
rect 13368 44552 13373 44608
rect 14043 44572 14048 44628
rect 14104 44572 14109 44628
rect 14043 44567 14109 44572
rect 14779 44628 14845 44633
rect 14779 44572 14784 44628
rect 14840 44572 14845 44628
rect 15518 44613 15578 44748
rect 16246 44708 16252 44772
rect 16316 44708 16322 44772
rect 16982 44728 16988 44792
rect 17052 44728 17058 44792
rect 24342 44749 24348 44813
rect 24412 44749 24418 44813
rect 16254 44613 16314 44708
rect 14779 44567 14845 44572
rect 15515 44608 15581 44613
rect 13307 44547 13373 44552
rect 15515 44552 15520 44608
rect 15576 44552 15581 44608
rect 15515 44547 15581 44552
rect 16251 44608 16317 44613
rect 16251 44552 16256 44608
rect 16312 44552 16317 44608
rect 16990 44573 17050 44728
rect 24350 44662 24410 44749
rect 24347 44657 24413 44662
rect 24347 44601 24352 44657
rect 24408 44601 24413 44657
rect 24347 44596 24413 44601
rect 16251 44547 16317 44552
rect 16987 44568 17053 44573
rect 9747 44530 11162 44532
rect 9747 44527 9813 44530
rect 16987 44512 16992 44568
rect 17048 44512 17053 44568
rect 16987 44507 17053 44512
rect 30971 44404 31035 44410
rect 8294 44342 30971 44402
rect 6627 44150 6693 44153
rect 8068 44152 8132 44158
rect 6627 44148 8068 44150
rect 6627 44092 6632 44148
rect 6688 44092 8068 44148
rect 6627 44090 8068 44092
rect 6627 44087 6693 44090
rect 8294 44145 8354 44342
rect 30971 44334 31035 44340
rect 8068 44082 8132 44088
rect 8289 44140 8359 44145
rect 8289 44080 8294 44140
rect 8354 44080 8359 44140
rect 22401 44086 22465 44092
rect 8289 44075 8359 44080
rect 20899 44024 22401 44084
rect 3147 43730 3213 43733
rect 3147 43728 3650 43730
rect 3147 43672 3152 43728
rect 3208 43672 3650 43728
rect 3147 43670 3650 43672
rect 3147 43667 3213 43670
rect 3590 42630 3650 43670
rect 9345 43650 9415 43655
rect 9345 43590 9350 43650
rect 9410 43590 9415 43650
rect 9345 43585 9415 43590
rect 9350 43418 9410 43585
rect 9348 43412 9412 43418
rect 9348 43342 9412 43348
rect 11564 43223 11570 43287
rect 11634 43285 11640 43287
rect 20899 43285 20959 44024
rect 22401 44016 22465 44022
rect 22413 43926 22477 43932
rect 11634 43225 20959 43285
rect 21071 43864 22413 43924
rect 11634 43223 11640 43225
rect 11732 43010 11738 43074
rect 11802 43072 11808 43074
rect 21071 43072 21131 43864
rect 22413 43856 22477 43862
rect 21278 43755 21342 43761
rect 22405 43755 22469 43761
rect 21342 43693 22405 43753
rect 21278 43685 21342 43691
rect 22405 43685 22469 43691
rect 22392 43545 22456 43551
rect 21438 43481 21444 43545
rect 21508 43543 21514 43545
rect 21508 43483 22392 43543
rect 21508 43481 21514 43483
rect 22392 43475 22456 43481
rect 22387 43291 22451 43297
rect 21615 43227 21621 43291
rect 21685 43289 21691 43291
rect 21685 43229 22387 43289
rect 21685 43227 21691 43229
rect 22387 43221 22451 43227
rect 11802 43012 21131 43072
rect 22393 43061 22457 43067
rect 11802 43010 11808 43012
rect 21796 42997 21802 43061
rect 21866 43059 21872 43061
rect 21866 42999 22393 43059
rect 21866 42997 21872 42999
rect 22393 42991 22457 42997
rect 10383 42901 10507 42913
rect 22404 42901 22499 42906
rect 10383 42900 22500 42901
rect 10383 42805 22404 42900
rect 22499 42805 22500 42900
rect 10383 42804 22500 42805
rect 10383 42716 10511 42804
rect 22404 42799 22499 42804
rect 9125 42630 9195 42635
rect 3590 42570 9130 42630
rect 9190 42570 9195 42630
rect 9125 42565 9195 42570
rect 9285 42410 9355 42415
rect 9150 42350 9290 42410
rect 9350 42350 9355 42410
rect 9285 42345 9355 42350
rect 1222 41730 1228 41732
rect 1090 41670 1228 41730
rect 1222 41668 1228 41670
rect 1292 41668 1298 41732
rect 982 39948 988 40012
rect 1052 39948 1058 40012
rect 990 39650 1050 39948
rect 9365 39010 9435 39015
rect 9270 38950 9370 39010
rect 9430 38950 9435 39010
rect 9365 38945 9435 38950
rect 945 37670 1015 37675
rect 770 37610 950 37670
rect 1010 37610 1015 37670
rect 945 37605 1015 37610
rect 10383 37008 10507 42716
rect 11370 42664 11440 42669
rect 11370 42604 11375 42664
rect 11435 42604 11440 42664
rect 11370 42599 11440 42604
rect 11375 42448 11435 42599
rect 11373 42442 11437 42448
rect 11373 42372 11437 42378
rect 12077 38161 12143 38164
rect 12412 38163 12476 38169
rect 12077 38159 12412 38161
rect 12077 38103 12082 38159
rect 12138 38103 12412 38159
rect 12077 38101 12412 38103
rect 12077 38098 12143 38101
rect 12412 38093 12476 38099
rect 12360 37520 12880 37540
rect 12360 37460 12380 37520
rect 12440 37460 12880 37520
rect 12360 37440 12880 37460
rect 9631 36888 10507 37008
rect 10383 36886 10507 36888
rect 1125 36290 1195 36295
rect 870 36230 1130 36290
rect 1190 36230 1195 36290
rect 1125 36225 1195 36230
rect 9425 34930 9495 34935
rect 9310 34870 9430 34930
rect 9490 34870 9495 34930
rect 9425 34865 9495 34870
rect 9342 34628 9348 34692
rect 9412 34628 9418 34692
rect 765 34270 835 34275
rect 765 34210 770 34270
rect 830 34210 990 34270
rect 765 34205 835 34210
rect 9350 33993 9410 34628
rect 9347 33988 9413 33993
rect 9347 33932 9352 33988
rect 9408 33932 9413 33988
rect 9347 33927 9413 33932
rect 5467 33190 5533 33193
rect 390 33188 5533 33190
rect 390 33132 5472 33188
rect 5528 33132 5533 33188
rect 390 33130 5533 33132
rect 5467 33127 5533 33130
rect 11885 32087 11951 32090
rect 12249 32089 12313 32095
rect 11885 32085 12249 32087
rect 11885 32029 11890 32085
rect 11946 32029 12249 32085
rect 11885 32027 12249 32029
rect 11885 32024 11951 32027
rect 12249 32019 12313 32025
rect 12360 31520 12780 31540
rect 12360 31460 12380 31520
rect 12440 31460 12780 31520
rect 12360 31440 12780 31460
rect 11685 26057 11751 26060
rect 12085 26059 12149 26065
rect 11685 26055 12085 26057
rect 11685 25999 11690 26055
rect 11746 25999 12085 26055
rect 11685 25997 12085 25999
rect 11685 25994 11751 25997
rect 12085 25989 12149 25995
rect 12360 25520 12840 25540
rect 12360 25460 12380 25520
rect 12440 25460 12840 25520
rect 12360 25440 12840 25460
rect 11562 20101 11628 20104
rect 11925 20103 11989 20109
rect 11562 20099 11925 20101
rect 11562 20043 11567 20099
rect 11623 20043 11925 20099
rect 11562 20041 11925 20043
rect 11562 20038 11628 20041
rect 11925 20033 11989 20039
rect 12360 19520 12840 19540
rect 12360 19460 12380 19520
rect 12440 19460 12840 19520
rect 12360 19440 12840 19460
rect 11732 14119 11738 14183
rect 11802 14119 11808 14183
rect 11740 14054 11800 14119
rect 11737 14049 11803 14054
rect 11737 13993 11742 14049
rect 11798 13993 11803 14049
rect 11737 13988 11803 13993
rect 12360 13520 12820 13540
rect 12360 13460 12380 13520
rect 12440 13460 12820 13520
rect 12360 13440 12820 13460
rect 11564 8249 11570 8313
rect 11634 8249 11640 8313
rect 11572 8135 11632 8249
rect 11569 8130 11635 8135
rect 11569 8074 11574 8130
rect 11630 8074 11635 8130
rect 11569 8069 11635 8074
rect 12360 7520 12820 7540
rect 12360 7460 12380 7520
rect 12440 7460 12820 7520
rect 12360 7440 12820 7460
rect 11367 2413 11373 2477
rect 11437 2413 11443 2477
rect 11375 2238 11435 2413
rect 11372 2233 11438 2238
rect 11372 2177 11377 2233
rect 11433 2177 11438 2233
rect 11372 2172 11438 2177
rect 12360 1520 12800 1540
rect 12360 1460 12380 1520
rect 12440 1460 12800 1520
rect 12360 1440 12800 1460
rect 30510 829 31462 830
rect 30510 825 31283 829
rect 30510 655 30515 825
rect 30685 655 31283 825
rect 30510 651 31283 655
rect 31461 651 31467 829
rect 30510 650 31462 651
<< via3 >>
rect 8156 44688 8220 44752
rect 10364 44708 10428 44772
rect 11100 44728 11164 44792
rect 11836 44728 11900 44792
rect 12572 44748 12636 44812
rect 13308 44748 13372 44812
rect 14044 44748 14108 44812
rect 988 44528 1052 44592
rect 14780 44728 14844 44792
rect 15516 44748 15580 44812
rect 16252 44708 16316 44772
rect 16988 44728 17052 44792
rect 24348 44749 24412 44813
rect 8068 44088 8132 44152
rect 30971 44340 31035 44404
rect 9348 43348 9412 43412
rect 11570 43223 11634 43287
rect 22401 44022 22465 44086
rect 11738 43010 11802 43074
rect 22413 43862 22477 43926
rect 21278 43691 21342 43755
rect 22405 43691 22469 43755
rect 21444 43481 21508 43545
rect 22392 43481 22456 43545
rect 21621 43227 21685 43291
rect 22387 43227 22451 43291
rect 21802 42997 21866 43061
rect 22393 42997 22457 43061
rect 22404 42805 22499 42900
rect 1228 41668 1292 41732
rect 988 39948 1052 40012
rect 11373 42378 11437 42442
rect 12412 38099 12476 38163
rect 9348 34628 9412 34692
rect 12249 32025 12313 32089
rect 12085 25995 12149 26059
rect 11925 20039 11989 20103
rect 11738 14119 11802 14183
rect 11570 8249 11634 8313
rect 11373 2413 11437 2477
rect 31283 651 31461 829
<< metal4 >>
rect 798 44773 858 45152
rect 1534 44773 1594 45152
rect 2270 44773 2330 45152
rect 3006 44773 3066 45152
rect 3742 44773 3802 45152
rect 4478 44773 4538 45152
rect 5214 44773 5274 45152
rect 5950 44773 6010 45152
rect 798 44713 6010 44773
rect 200 44050 500 44152
rect 798 44050 858 44713
rect 987 44592 1053 44593
rect 987 44528 988 44592
rect 1052 44590 1053 44592
rect 6686 44590 6746 45152
rect 1052 44530 6746 44590
rect 1052 44528 1053 44530
rect 987 44527 1053 44528
rect 7422 44430 7482 45152
rect 8158 44753 8218 45152
rect 8155 44752 8221 44753
rect 8155 44688 8156 44752
rect 8220 44688 8221 44752
rect 8155 44687 8221 44688
rect 200 43990 858 44050
rect 990 44370 7482 44430
rect 200 34800 500 43990
rect 990 40013 1050 44370
rect 8067 44152 8133 44153
rect 8067 44088 8068 44152
rect 8132 44150 8133 44152
rect 8894 44150 8954 45152
rect 8132 44090 8954 44150
rect 8132 44088 8133 44090
rect 8067 44087 8133 44088
rect 9630 43890 9690 45152
rect 10366 44773 10426 45152
rect 11102 44793 11162 45152
rect 11838 44793 11898 45152
rect 12574 44813 12634 45152
rect 13310 44813 13370 45152
rect 14046 44813 14106 45152
rect 12571 44812 12637 44813
rect 11099 44792 11165 44793
rect 10363 44772 10429 44773
rect 10363 44708 10364 44772
rect 10428 44708 10429 44772
rect 11099 44728 11100 44792
rect 11164 44728 11165 44792
rect 11099 44727 11165 44728
rect 11835 44792 11901 44793
rect 11835 44728 11836 44792
rect 11900 44728 11901 44792
rect 12571 44748 12572 44812
rect 12636 44748 12637 44812
rect 12571 44747 12637 44748
rect 13307 44812 13373 44813
rect 13307 44748 13308 44812
rect 13372 44748 13373 44812
rect 13307 44747 13373 44748
rect 14043 44812 14109 44813
rect 14043 44748 14044 44812
rect 14108 44748 14109 44812
rect 14782 44793 14842 45152
rect 15518 44813 15578 45152
rect 15515 44812 15581 44813
rect 14043 44747 14109 44748
rect 14779 44792 14845 44793
rect 11835 44727 11901 44728
rect 14779 44728 14780 44792
rect 14844 44728 14845 44792
rect 15515 44748 15516 44812
rect 15580 44748 15581 44812
rect 16254 44773 16314 45152
rect 16990 44793 17050 45152
rect 16987 44792 17053 44793
rect 15515 44747 15581 44748
rect 16251 44772 16317 44773
rect 14779 44727 14845 44728
rect 10363 44707 10429 44708
rect 16251 44708 16252 44772
rect 16316 44708 16317 44772
rect 16987 44728 16988 44792
rect 17052 44728 17053 44792
rect 16987 44727 17053 44728
rect 16251 44707 16317 44708
rect 17726 44200 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44814 24410 45152
rect 24347 44813 24413 44814
rect 24347 44749 24348 44813
rect 24412 44749 24413 44813
rect 24347 44748 24413 44749
rect 1230 43830 9690 43890
rect 9800 43853 22293 44200
rect 22400 44086 22466 44087
rect 22400 44022 22401 44086
rect 22465 44084 22466 44086
rect 25086 44084 25146 45152
rect 22465 44024 25146 44084
rect 22465 44022 22466 44024
rect 22400 44021 22466 44022
rect 22412 43926 22478 43927
rect 22412 43862 22413 43926
rect 22477 43924 22478 43926
rect 25822 43924 25882 45152
rect 22477 43864 25882 43924
rect 22477 43862 22478 43864
rect 22412 43861 22478 43862
rect 1230 41733 1290 43830
rect 9800 43600 10122 43853
rect 21277 43755 21343 43756
rect 21277 43691 21278 43755
rect 21342 43691 21343 43755
rect 21277 43690 21343 43691
rect 9347 43412 9413 43413
rect 9347 43348 9348 43412
rect 9412 43348 9413 43412
rect 9347 43347 9413 43348
rect 1227 41732 1293 41733
rect 1227 41668 1228 41732
rect 1292 41668 1293 41732
rect 1227 41667 1293 41668
rect 987 40012 1053 40013
rect 987 39948 988 40012
rect 1052 39948 1053 40012
rect 987 39947 1053 39948
rect 2400 34800 2700 35100
rect 200 34500 2700 34800
rect 8293 34505 8570 35267
rect 9350 34693 9410 43347
rect 9347 34692 9413 34693
rect 9347 34628 9348 34692
rect 9412 34628 9413 34692
rect 9347 34627 9413 34628
rect 9800 34505 10100 43600
rect 21280 43471 21340 43690
rect 21443 43545 21509 43546
rect 21443 43481 21444 43545
rect 21508 43481 21509 43545
rect 21443 43480 21509 43481
rect 11927 43411 21340 43471
rect 11569 43287 11635 43288
rect 11569 43223 11570 43287
rect 11634 43223 11635 43287
rect 11569 43222 11635 43223
rect 11372 42442 11438 42443
rect 11372 42378 11373 42442
rect 11437 42378 11438 42442
rect 11372 42377 11438 42378
rect 200 1000 500 34500
rect 8293 34187 10100 34505
rect 9800 894 10100 34187
rect 11375 2478 11435 42377
rect 11572 8314 11632 43222
rect 11737 43074 11803 43075
rect 11737 43010 11738 43074
rect 11802 43010 11803 43074
rect 11737 43009 11803 43010
rect 11740 14184 11800 43009
rect 11927 20104 11987 43411
rect 21446 43279 21506 43480
rect 12087 43219 21506 43279
rect 21620 43291 21686 43292
rect 21620 43227 21621 43291
rect 21685 43227 21686 43291
rect 21620 43226 21686 43227
rect 12087 26060 12147 43219
rect 21623 43071 21683 43226
rect 12251 43011 21683 43071
rect 21801 43061 21867 43062
rect 12251 32090 12311 43011
rect 21801 42997 21802 43061
rect 21866 42997 21867 43061
rect 21801 42996 21867 42997
rect 21804 42878 21864 42996
rect 12411 42818 21864 42878
rect 12411 42753 12543 42818
rect 12411 42752 12474 42753
rect 12414 38164 12474 42752
rect 12411 38163 12477 38164
rect 12411 38099 12412 38163
rect 12476 38099 12477 38163
rect 12411 38098 12477 38099
rect 12248 32089 12314 32090
rect 12248 32025 12249 32089
rect 12313 32025 12314 32089
rect 12248 32024 12314 32025
rect 12084 26059 12150 26060
rect 12084 25995 12085 26059
rect 12149 25995 12150 26059
rect 12084 25994 12150 25995
rect 11924 20103 11990 20104
rect 11924 20039 11925 20103
rect 11989 20039 11990 20103
rect 11924 20038 11990 20039
rect 11737 14183 11803 14184
rect 11737 14119 11738 14183
rect 11802 14119 11803 14183
rect 11737 14118 11803 14119
rect 11569 8313 11635 8314
rect 11569 8249 11570 8313
rect 11634 8249 11635 8313
rect 11569 8248 11635 8249
rect 11372 2477 11438 2478
rect 11372 2413 11373 2477
rect 11437 2413 11438 2477
rect 11372 2412 11438 2413
rect 15650 894 15950 42546
rect 21946 1559 22293 43853
rect 22404 43755 22470 43756
rect 22404 43691 22405 43755
rect 22469 43753 22470 43755
rect 26558 43753 26618 45152
rect 22469 43693 26618 43753
rect 22469 43691 22470 43693
rect 22404 43690 22470 43691
rect 22391 43545 22457 43546
rect 22391 43481 22392 43545
rect 22456 43543 22457 43545
rect 27294 43543 27354 45152
rect 22456 43483 27354 43543
rect 22456 43481 22457 43483
rect 22391 43480 22457 43481
rect 22386 43291 22452 43292
rect 22386 43227 22387 43291
rect 22451 43289 22452 43291
rect 28030 43289 28090 45152
rect 22451 43229 28090 43289
rect 22451 43227 22452 43229
rect 22386 43226 22452 43227
rect 22392 43061 22458 43062
rect 22392 42997 22393 43061
rect 22457 43059 22458 43061
rect 28766 43059 28826 45152
rect 29502 44952 29562 45152
rect 30238 45087 30298 45152
rect 30173 44952 30298 45087
rect 30974 44999 31034 45152
rect 30973 44952 31034 44999
rect 31710 44952 31770 45152
rect 30173 43059 30297 44952
rect 30973 44405 31033 44952
rect 30970 44404 31036 44405
rect 30970 44340 30971 44404
rect 31035 44340 31036 44404
rect 30970 44339 31036 44340
rect 22457 42999 28826 43059
rect 22457 42997 22458 42999
rect 22392 42996 22458 42997
rect 30187 42901 30284 43059
rect 22403 42900 30284 42901
rect 22403 42805 22404 42900
rect 22499 42805 30284 42900
rect 22403 42804 30284 42805
rect 28857 894 29157 42560
rect 9800 594 29157 894
rect 31282 829 31462 830
rect 31282 651 31283 829
rect 31461 651 31462 829
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 651
use psu_sequencer  psu_sequencer_0 ~/projects/adia/adia_psu_full_test/mag
timestamp 1717221846
transform 1 0 550 0 1 32800
box 0 0 9204 11348
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_0
timestamp 1717221846
transform 1 0 4166 0 1 19020
box -1786 -1640 1786 1640
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_0
timestamp 1717221846
transform 1 0 22398 0 1 3840
box -9798 -2840 9798 2840
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_1
timestamp 1717221846
transform 1 0 22398 0 1 39840
box -9798 -2840 9798 2840
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_2
timestamp 1717221846
transform 1 0 22398 0 1 33840
box -9798 -2840 9798 2840
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_3
timestamp 1717221846
transform 1 0 22398 0 1 27840
box -9798 -2840 9798 2840
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_4
timestamp 1717221846
transform 1 0 22398 0 1 21840
box -9798 -2840 9798 2840
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_5
timestamp 1717221846
transform 1 0 22398 0 1 15840
box -9798 -2840 9798 2840
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_6
timestamp 1717221846
transform 1 0 22398 0 1 9840
box -9798 -2840 9798 2840
use sky130_fd_pr__nfet_01v8_EDB9KC  sky130_fd_pr__nfet_01v8_EDB9KC_0
timestamp 1717221846
transform 1 0 4115 0 1 22256
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_0
timestamp 1717221846
transform 1 0 2531 0 1 23292
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_1
timestamp 1717221846
transform 0 1 12118 -1 0 7693
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_2
timestamp 1717221846
transform 0 1 12118 -1 0 1693
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_3
timestamp 1717221846
transform 0 1 12118 -1 0 19693
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_4
timestamp 1717221846
transform 0 1 12118 -1 0 13693
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_5
timestamp 1717221846
transform 0 1 12118 -1 0 31693
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_6
timestamp 1717221846
transform 0 1 12118 -1 0 25693
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_7
timestamp 1717221846
transform 0 1 12118 -1 0 37693
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_0
timestamp 1717221846
transform 1 0 2993 0 1 23293
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_1
timestamp 1717221846
transform 0 1 12119 -1 0 7231
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_2
timestamp 1717221846
transform 0 1 12119 -1 0 1231
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_3
timestamp 1717221846
transform 0 1 12119 -1 0 19231
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_4
timestamp 1717221846
transform 0 1 12119 -1 0 13231
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_5
timestamp 1717221846
transform 0 1 12119 -1 0 31231
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_6
timestamp 1717221846
transform 0 1 12119 -1 0 25231
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_7
timestamp 1717221846
transform 0 1 12119 -1 0 37231
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_UAQRRG  sky130_fd_pr__pfet_01v8_UAQRRG_0
timestamp 1717221846
transform 1 0 3203 0 1 21977
box -211 -319 211 319
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 11398 0 -1 7592
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1717221846
transform 1 0 11398 0 -1 1592
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1717221846
transform 1 0 11398 0 -1 13592
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1717221846
transform -1 0 1934 0 -1 22992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1717221846
transform 1 0 11398 0 -1 31592
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1717221846
transform 1 0 11398 0 -1 25592
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1717221846
transform 1 0 11398 0 -1 37592
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_7
timestamp 1717221846
transform 1 0 11398 0 -1 19592
box -38 -48 314 592
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
