magic
tech sky130A
magscale 1 2
timestamp 1717221846
<< viali >>
rect 2973 8585 3007 8619
rect 6561 8585 6595 8619
rect 7113 8585 7147 8619
rect 7573 8585 7607 8619
rect 2421 8517 2455 8551
rect 4721 8517 4755 8551
rect 4813 8517 4847 8551
rect 1777 8449 1811 8483
rect 2053 8449 2087 8483
rect 3065 8449 3099 8483
rect 3433 8449 3467 8483
rect 3617 8449 3651 8483
rect 4353 8449 4387 8483
rect 4537 8449 4571 8483
rect 4905 8449 4939 8483
rect 5365 8449 5399 8483
rect 6469 8449 6503 8483
rect 6929 8449 6963 8483
rect 7665 8449 7699 8483
rect 4077 8381 4111 8415
rect 5549 8381 5583 8415
rect 1501 8313 1535 8347
rect 5089 8313 5123 8347
rect 3249 8245 3283 8279
rect 5181 8245 5215 8279
rect 1501 8041 1535 8075
rect 1961 8041 1995 8075
rect 4997 8041 5031 8075
rect 6837 8041 6871 8075
rect 3065 7973 3099 8007
rect 2145 7837 2179 7871
rect 2421 7837 2455 7871
rect 2605 7837 2639 7871
rect 2789 7837 2823 7871
rect 4353 7837 4387 7871
rect 6745 7837 6779 7871
rect 7021 7837 7055 7871
rect 7389 7837 7423 7871
rect 7481 7837 7515 7871
rect 1777 7769 1811 7803
rect 2513 7769 2547 7803
rect 3249 7769 3283 7803
rect 6469 7769 6503 7803
rect 7113 7769 7147 7803
rect 7205 7769 7239 7803
rect 2237 7701 2271 7735
rect 3801 7701 3835 7735
rect 7665 7701 7699 7735
rect 1685 7497 1719 7531
rect 2329 7497 2363 7531
rect 6101 7497 6135 7531
rect 7113 7497 7147 7531
rect 2053 7429 2087 7463
rect 1409 7361 1443 7395
rect 1869 7361 1903 7395
rect 2145 7361 2179 7395
rect 4077 7361 4111 7395
rect 4445 7361 4479 7395
rect 5273 7361 5307 7395
rect 6929 7361 6963 7395
rect 7297 7361 7331 7395
rect 7389 7361 7423 7395
rect 7481 7361 7515 7395
rect 7665 7361 7699 7395
rect 3801 7293 3835 7327
rect 4721 7293 4755 7327
rect 5457 7293 5491 7327
rect 4629 7225 4663 7259
rect 1593 7157 1627 7191
rect 6377 7157 6411 7191
rect 5641 6953 5675 6987
rect 1685 6885 1719 6919
rect 3249 6817 3283 6851
rect 7389 6817 7423 6851
rect 1501 6749 1535 6783
rect 2533 6749 2567 6783
rect 2789 6749 2823 6783
rect 2881 6749 2915 6783
rect 3985 6749 4019 6783
rect 4261 6749 4295 6783
rect 5457 6749 5491 6783
rect 2329 6681 2363 6715
rect 2697 6681 2731 6715
rect 3525 6681 3559 6715
rect 3801 6681 3835 6715
rect 7113 6681 7147 6715
rect 2237 6613 2271 6647
rect 3065 6613 3099 6647
rect 4169 6613 4203 6647
rect 5273 6613 5307 6647
rect 1409 6409 1443 6443
rect 3663 6409 3697 6443
rect 6561 6341 6595 6375
rect 7389 6341 7423 6375
rect 1593 6273 1627 6307
rect 1685 6273 1719 6307
rect 5825 6273 5859 6307
rect 6377 6273 6411 6307
rect 6653 6273 6687 6307
rect 6745 6273 6779 6307
rect 7205 6273 7239 6307
rect 7297 6273 7331 6307
rect 7573 6273 7607 6307
rect 1869 6205 1903 6239
rect 2237 6205 2271 6239
rect 3801 6205 3835 6239
rect 4077 6205 4111 6239
rect 6929 6137 6963 6171
rect 5549 6069 5583 6103
rect 6101 6069 6135 6103
rect 7021 6069 7055 6103
rect 4445 5865 4479 5899
rect 5365 5865 5399 5899
rect 7665 5865 7699 5899
rect 5641 5729 5675 5763
rect 2053 5661 2087 5695
rect 2237 5661 2271 5695
rect 2421 5661 2455 5695
rect 2697 5637 2731 5671
rect 3065 5661 3099 5695
rect 3157 5661 3191 5695
rect 3249 5661 3283 5695
rect 3433 5661 3467 5695
rect 3893 5661 3927 5695
rect 4997 5661 5031 5695
rect 5181 5661 5215 5695
rect 7481 5661 7515 5695
rect 2145 5593 2179 5627
rect 4261 5593 4295 5627
rect 5917 5593 5951 5627
rect 1869 5525 1903 5559
rect 2513 5525 2547 5559
rect 2881 5525 2915 5559
rect 7389 5525 7423 5559
rect 6469 5321 6503 5355
rect 6837 5321 6871 5355
rect 1777 5253 1811 5287
rect 2605 5253 2639 5287
rect 6193 5253 6227 5287
rect 1961 5185 1995 5219
rect 2397 5185 2431 5219
rect 2513 5185 2547 5219
rect 2789 5185 2823 5219
rect 2973 5185 3007 5219
rect 3893 5185 3927 5219
rect 6653 5185 6687 5219
rect 7389 5185 7423 5219
rect 7757 5185 7791 5219
rect 3985 5117 4019 5151
rect 4077 5117 4111 5151
rect 3157 5049 3191 5083
rect 1501 4981 1535 5015
rect 2145 4981 2179 5015
rect 2237 4981 2271 5015
rect 3525 4981 3559 5015
rect 4721 4981 4755 5015
rect 7573 4981 7607 5015
rect 4537 4777 4571 4811
rect 6745 4777 6779 4811
rect 2605 4709 2639 4743
rect 3433 4641 3467 4675
rect 3985 4641 4019 4675
rect 7665 4641 7699 4675
rect 1777 4573 1811 4607
rect 2329 4573 2363 4607
rect 2789 4573 2823 4607
rect 4169 4573 4203 4607
rect 5273 4573 5307 4607
rect 1409 4505 1443 4539
rect 1961 4505 1995 4539
rect 4077 4505 4111 4539
rect 4813 4505 4847 4539
rect 5181 4505 5215 4539
rect 2881 4437 2915 4471
rect 3249 4437 3283 4471
rect 3341 4437 3375 4471
rect 7113 4437 7147 4471
rect 6101 4233 6135 4267
rect 6377 4233 6411 4267
rect 7757 4233 7791 4267
rect 4629 4165 4663 4199
rect 7389 4165 7423 4199
rect 1869 4097 1903 4131
rect 1961 4097 1995 4131
rect 2145 4097 2179 4131
rect 4353 4097 4387 4131
rect 6929 4097 6963 4131
rect 7205 4097 7239 4131
rect 7481 4097 7515 4131
rect 7573 4097 7607 4131
rect 2421 4029 2455 4063
rect 2789 4029 2823 4063
rect 2329 3893 2363 3927
rect 4215 3893 4249 3927
rect 7665 3689 7699 3723
rect 1869 3553 1903 3587
rect 5825 3553 5859 3587
rect 5917 3553 5951 3587
rect 3801 3485 3835 3519
rect 2145 3417 2179 3451
rect 5549 3417 5583 3451
rect 6193 3417 6227 3451
rect 3617 3349 3651 3383
rect 3985 3349 4019 3383
rect 4077 3349 4111 3383
rect 2145 3145 2179 3179
rect 2513 3145 2547 3179
rect 4445 3145 4479 3179
rect 4813 3145 4847 3179
rect 5917 3145 5951 3179
rect 7113 3145 7147 3179
rect 4353 3077 4387 3111
rect 6561 3077 6595 3111
rect 1869 3009 1903 3043
rect 2053 3009 2087 3043
rect 2329 3009 2363 3043
rect 5273 3009 5307 3043
rect 6745 3009 6779 3043
rect 7021 3009 7055 3043
rect 7297 3009 7331 3043
rect 7389 3009 7423 3043
rect 7481 3009 7515 3043
rect 7665 3009 7699 3043
rect 2605 2941 2639 2975
rect 4905 2941 4939 2975
rect 4997 2941 5031 2975
rect 6929 2941 6963 2975
rect 1777 2805 1811 2839
rect 3801 2601 3835 2635
rect 3617 2533 3651 2567
rect 1869 2465 1903 2499
rect 4169 2465 4203 2499
rect 5733 2465 5767 2499
rect 3985 2397 4019 2431
rect 4353 2397 4387 2431
rect 4813 2397 4847 2431
rect 5181 2397 5215 2431
rect 5609 2397 5643 2431
rect 5825 2397 5859 2431
rect 6837 2397 6871 2431
rect 7021 2397 7055 2431
rect 2145 2329 2179 2363
rect 4721 2329 4755 2363
rect 6469 2329 6503 2363
rect 5365 2261 5399 2295
rect 7113 2261 7147 2295
<< metal1 >>
rect 2774 8848 2780 8900
rect 2832 8888 2838 8900
rect 2958 8888 2964 8900
rect 2832 8860 2964 8888
rect 2832 8848 2838 8860
rect 2958 8848 2964 8860
rect 3016 8848 3022 8900
rect 4614 8780 4620 8832
rect 4672 8820 4678 8832
rect 5258 8820 5264 8832
rect 4672 8792 5264 8820
rect 4672 8780 4678 8792
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 1104 8730 8096 8752
rect 1104 8678 2483 8730
rect 2535 8678 2547 8730
rect 2599 8678 2611 8730
rect 2663 8678 2675 8730
rect 2727 8678 2739 8730
rect 2791 8678 4230 8730
rect 4282 8678 4294 8730
rect 4346 8678 4358 8730
rect 4410 8678 4422 8730
rect 4474 8678 4486 8730
rect 4538 8678 5977 8730
rect 6029 8678 6041 8730
rect 6093 8678 6105 8730
rect 6157 8678 6169 8730
rect 6221 8678 6233 8730
rect 6285 8678 7724 8730
rect 7776 8678 7788 8730
rect 7840 8678 7852 8730
rect 7904 8678 7916 8730
rect 7968 8678 7980 8730
rect 8032 8678 8096 8730
rect 1104 8656 8096 8678
rect 2958 8576 2964 8628
rect 3016 8576 3022 8628
rect 3970 8616 3976 8628
rect 3620 8588 3976 8616
rect 2409 8551 2467 8557
rect 2409 8517 2421 8551
rect 2455 8548 2467 8551
rect 2866 8548 2872 8560
rect 2455 8520 2872 8548
rect 2455 8517 2467 8520
rect 2409 8511 2467 8517
rect 2866 8508 2872 8520
rect 2924 8508 2930 8560
rect 1670 8440 1676 8492
rect 1728 8480 1734 8492
rect 1765 8483 1823 8489
rect 1765 8480 1777 8483
rect 1728 8452 1777 8480
rect 1728 8440 1734 8452
rect 1765 8449 1777 8452
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 2222 8480 2228 8492
rect 2087 8452 2228 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 3050 8440 3056 8492
rect 3108 8440 3114 8492
rect 3620 8489 3648 8588
rect 3970 8576 3976 8588
rect 4028 8616 4034 8628
rect 5534 8616 5540 8628
rect 4028 8588 5540 8616
rect 4028 8576 4034 8588
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 5868 8588 6561 8616
rect 5868 8576 5874 8588
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 6549 8579 6607 8585
rect 7098 8576 7104 8628
rect 7156 8576 7162 8628
rect 7561 8619 7619 8625
rect 7561 8585 7573 8619
rect 7607 8616 7619 8619
rect 9030 8616 9036 8628
rect 7607 8588 9036 8616
rect 7607 8585 7619 8588
rect 7561 8579 7619 8585
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 4709 8551 4767 8557
rect 4709 8548 4721 8551
rect 4172 8520 4721 8548
rect 4172 8492 4200 8520
rect 4709 8517 4721 8520
rect 4755 8517 4767 8551
rect 4709 8511 4767 8517
rect 4801 8551 4859 8557
rect 4801 8517 4813 8551
rect 4847 8548 4859 8551
rect 4847 8520 5120 8548
rect 4847 8517 4859 8520
rect 4801 8511 4859 8517
rect 5092 8492 5120 8520
rect 5258 8508 5264 8560
rect 5316 8548 5322 8560
rect 6362 8548 6368 8560
rect 5316 8520 6368 8548
rect 5316 8508 5322 8520
rect 6362 8508 6368 8520
rect 6420 8508 6426 8560
rect 3421 8483 3479 8489
rect 3421 8480 3433 8483
rect 3160 8452 3433 8480
rect 3160 8356 3188 8452
rect 3421 8449 3433 8452
rect 3467 8449 3479 8483
rect 3421 8443 3479 8449
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 4154 8440 4160 8492
rect 4212 8440 4218 8492
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 4614 8480 4620 8492
rect 4571 8452 4620 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 3878 8372 3884 8424
rect 3936 8412 3942 8424
rect 4065 8415 4123 8421
rect 4065 8412 4077 8415
rect 3936 8384 4077 8412
rect 3936 8372 3942 8384
rect 4065 8381 4077 8384
rect 4111 8381 4123 8415
rect 4356 8412 4384 8443
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 4893 8483 4951 8489
rect 4893 8449 4905 8483
rect 4939 8480 4951 8483
rect 4982 8480 4988 8492
rect 4939 8452 4988 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 5074 8440 5080 8492
rect 5132 8440 5138 8492
rect 5276 8480 5304 8508
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 5276 8452 5365 8480
rect 5353 8449 5365 8452
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 5460 8452 5672 8480
rect 5460 8412 5488 8452
rect 4356 8384 5488 8412
rect 4065 8375 4123 8381
rect 5534 8372 5540 8424
rect 5592 8372 5598 8424
rect 5644 8412 5672 8452
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 6457 8483 6515 8489
rect 6457 8480 6469 8483
rect 5776 8452 6469 8480
rect 5776 8440 5782 8452
rect 6457 8449 6469 8452
rect 6503 8449 6515 8483
rect 6457 8443 6515 8449
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 6880 8452 6929 8480
rect 6880 8440 6886 8452
rect 6917 8449 6929 8452
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 7616 8452 7665 8480
rect 7616 8440 7622 8452
rect 7653 8449 7665 8452
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 6546 8412 6552 8424
rect 5644 8384 6552 8412
rect 6546 8372 6552 8384
rect 6604 8372 6610 8424
rect 1489 8347 1547 8353
rect 1489 8313 1501 8347
rect 1535 8313 1547 8347
rect 1489 8307 1547 8313
rect 658 8236 664 8288
rect 716 8276 722 8288
rect 1504 8276 1532 8307
rect 3142 8304 3148 8356
rect 3200 8304 3206 8356
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8344 5135 8347
rect 6270 8344 6276 8356
rect 5123 8316 6276 8344
rect 5123 8313 5135 8316
rect 5077 8307 5135 8313
rect 6270 8304 6276 8316
rect 6328 8304 6334 8356
rect 716 8248 1532 8276
rect 716 8236 722 8248
rect 2498 8236 2504 8288
rect 2556 8276 2562 8288
rect 3237 8279 3295 8285
rect 3237 8276 3249 8279
rect 2556 8248 3249 8276
rect 2556 8236 2562 8248
rect 3237 8245 3249 8248
rect 3283 8245 3295 8279
rect 3237 8239 3295 8245
rect 5166 8236 5172 8288
rect 5224 8236 5230 8288
rect 1104 8186 8096 8208
rect 1104 8134 1823 8186
rect 1875 8134 1887 8186
rect 1939 8134 1951 8186
rect 2003 8134 2015 8186
rect 2067 8134 2079 8186
rect 2131 8134 3570 8186
rect 3622 8134 3634 8186
rect 3686 8134 3698 8186
rect 3750 8134 3762 8186
rect 3814 8134 3826 8186
rect 3878 8134 5317 8186
rect 5369 8134 5381 8186
rect 5433 8134 5445 8186
rect 5497 8134 5509 8186
rect 5561 8134 5573 8186
rect 5625 8134 7064 8186
rect 7116 8134 7128 8186
rect 7180 8134 7192 8186
rect 7244 8134 7256 8186
rect 7308 8134 7320 8186
rect 7372 8134 8096 8186
rect 1104 8112 8096 8134
rect 1486 8032 1492 8084
rect 1544 8032 1550 8084
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2222 8072 2228 8084
rect 1995 8044 2228 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 2406 8032 2412 8084
rect 2464 8072 2470 8084
rect 4985 8075 5043 8081
rect 4985 8072 4997 8075
rect 2464 8044 4997 8072
rect 2464 8032 2470 8044
rect 4985 8041 4997 8044
rect 5031 8041 5043 8075
rect 4985 8035 5043 8041
rect 3053 8007 3111 8013
rect 1504 7976 2728 8004
rect 1504 7812 1532 7976
rect 2498 7936 2504 7948
rect 2148 7908 2504 7936
rect 1670 7828 1676 7880
rect 1728 7828 1734 7880
rect 2148 7877 2176 7908
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 2700 7880 2728 7976
rect 3053 7973 3065 8007
rect 3099 8004 3111 8007
rect 4798 8004 4804 8016
rect 3099 7976 4804 8004
rect 3099 7973 3111 7976
rect 3053 7967 3111 7973
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 5000 7936 5028 8035
rect 6270 8032 6276 8084
rect 6328 8072 6334 8084
rect 6328 8044 6776 8072
rect 6328 8032 6334 8044
rect 6748 8004 6776 8044
rect 6822 8032 6828 8084
rect 6880 8032 6886 8084
rect 6748 7976 7512 8004
rect 6914 7936 6920 7948
rect 4080 7908 4660 7936
rect 5000 7908 6920 7936
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 2406 7868 2412 7880
rect 2280 7840 2412 7868
rect 2280 7828 2286 7840
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7864 2651 7871
rect 2682 7864 2688 7880
rect 2639 7837 2688 7864
rect 2593 7836 2688 7837
rect 2593 7831 2651 7836
rect 2682 7828 2688 7836
rect 2740 7828 2746 7880
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 4080 7868 4108 7908
rect 4632 7880 4660 7908
rect 6914 7896 6920 7908
rect 6972 7936 6978 7948
rect 6972 7908 7052 7936
rect 6972 7896 6978 7908
rect 2823 7840 4108 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 1486 7760 1492 7812
rect 1544 7760 1550 7812
rect 1688 7732 1716 7828
rect 1762 7760 1768 7812
rect 1820 7760 1826 7812
rect 2501 7803 2559 7809
rect 2501 7769 2513 7803
rect 2547 7800 2559 7803
rect 2866 7800 2872 7812
rect 2547 7772 2872 7800
rect 2547 7769 2559 7772
rect 2501 7763 2559 7769
rect 2866 7760 2872 7772
rect 2924 7760 2930 7812
rect 2225 7735 2283 7741
rect 2225 7732 2237 7735
rect 1688 7704 2237 7732
rect 2225 7701 2237 7704
rect 2271 7701 2283 7735
rect 2225 7695 2283 7701
rect 2314 7692 2320 7744
rect 2372 7732 2378 7744
rect 2976 7732 3004 7840
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4341 7871 4399 7877
rect 4341 7868 4353 7871
rect 4212 7840 4353 7868
rect 4212 7828 4218 7840
rect 4341 7837 4353 7840
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 4614 7828 4620 7880
rect 4672 7828 4678 7880
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 4764 7840 5382 7868
rect 4764 7828 4770 7840
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 7024 7877 7052 7908
rect 7484 7877 7512 7976
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 3237 7803 3295 7809
rect 3237 7769 3249 7803
rect 3283 7800 3295 7803
rect 3283 7772 5212 7800
rect 3283 7769 3295 7772
rect 3237 7763 3295 7769
rect 2372 7704 3004 7732
rect 2372 7692 2378 7704
rect 3326 7692 3332 7744
rect 3384 7732 3390 7744
rect 3789 7735 3847 7741
rect 3789 7732 3801 7735
rect 3384 7704 3801 7732
rect 3384 7692 3390 7704
rect 3789 7701 3801 7704
rect 3835 7701 3847 7735
rect 5184 7732 5212 7772
rect 6454 7760 6460 7812
rect 6512 7760 6518 7812
rect 7098 7760 7104 7812
rect 7156 7760 7162 7812
rect 7193 7803 7251 7809
rect 7193 7769 7205 7803
rect 7239 7769 7251 7803
rect 7392 7800 7420 7831
rect 8202 7828 8208 7880
rect 8260 7828 8266 7880
rect 8220 7800 8248 7828
rect 7392 7772 8248 7800
rect 7193 7763 7251 7769
rect 5534 7732 5540 7744
rect 5184 7704 5540 7732
rect 3789 7695 3847 7701
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 5810 7692 5816 7744
rect 5868 7732 5874 7744
rect 7208 7732 7236 7763
rect 5868 7704 7236 7732
rect 7653 7735 7711 7741
rect 5868 7692 5874 7704
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 8110 7732 8116 7744
rect 7699 7704 8116 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 1104 7642 8096 7664
rect 1104 7590 2483 7642
rect 2535 7590 2547 7642
rect 2599 7590 2611 7642
rect 2663 7590 2675 7642
rect 2727 7590 2739 7642
rect 2791 7590 4230 7642
rect 4282 7590 4294 7642
rect 4346 7590 4358 7642
rect 4410 7590 4422 7642
rect 4474 7590 4486 7642
rect 4538 7590 5977 7642
rect 6029 7590 6041 7642
rect 6093 7590 6105 7642
rect 6157 7590 6169 7642
rect 6221 7590 6233 7642
rect 6285 7590 7724 7642
rect 7776 7590 7788 7642
rect 7840 7590 7852 7642
rect 7904 7590 7916 7642
rect 7968 7590 7980 7642
rect 8032 7590 8096 7642
rect 1104 7568 8096 7590
rect 1673 7531 1731 7537
rect 1673 7497 1685 7531
rect 1719 7528 1731 7531
rect 1762 7528 1768 7540
rect 1719 7500 1768 7528
rect 1719 7497 1731 7500
rect 1673 7491 1731 7497
rect 1762 7488 1768 7500
rect 1820 7488 1826 7540
rect 2317 7531 2375 7537
rect 2317 7497 2329 7531
rect 2363 7528 2375 7531
rect 2406 7528 2412 7540
rect 2363 7500 2412 7528
rect 2363 7497 2375 7500
rect 2317 7491 2375 7497
rect 2406 7488 2412 7500
rect 2464 7528 2470 7540
rect 4154 7528 4160 7540
rect 2464 7500 4160 7528
rect 2464 7488 2470 7500
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 5166 7488 5172 7540
rect 5224 7488 5230 7540
rect 6089 7531 6147 7537
rect 6089 7497 6101 7531
rect 6135 7528 6147 7531
rect 6454 7528 6460 7540
rect 6135 7500 6460 7528
rect 6135 7497 6147 7500
rect 6089 7491 6147 7497
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 7101 7531 7159 7537
rect 7101 7528 7113 7531
rect 6604 7500 7113 7528
rect 6604 7488 6610 7500
rect 7101 7497 7113 7500
rect 7147 7497 7159 7531
rect 7101 7491 7159 7497
rect 2041 7463 2099 7469
rect 2041 7460 2053 7463
rect 1688 7432 2053 7460
rect 1688 7404 1716 7432
rect 2041 7429 2053 7432
rect 2087 7460 2099 7463
rect 3694 7460 3700 7472
rect 2087 7432 2544 7460
rect 3358 7432 3700 7460
rect 2087 7429 2099 7432
rect 2041 7423 2099 7429
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 1670 7352 1676 7404
rect 1728 7352 1734 7404
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 2314 7392 2320 7404
rect 2179 7364 2320 7392
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 1872 7324 1900 7355
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 2516 7392 2544 7432
rect 3694 7420 3700 7432
rect 3752 7460 3758 7472
rect 4706 7460 4712 7472
rect 3752 7432 4712 7460
rect 3752 7420 3758 7432
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 2516 7364 2636 7392
rect 2498 7324 2504 7336
rect 1872 7296 2504 7324
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 2608 7324 2636 7364
rect 4062 7352 4068 7404
rect 4120 7352 4126 7404
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 5184 7392 5212 7488
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 5592 7432 6592 7460
rect 5592 7420 5598 7432
rect 6564 7404 6592 7432
rect 6656 7432 7696 7460
rect 6656 7404 6684 7432
rect 4479 7364 5212 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 5810 7392 5816 7404
rect 5316 7364 5816 7392
rect 5316 7352 5322 7364
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 6362 7352 6368 7404
rect 6420 7352 6426 7404
rect 6546 7352 6552 7404
rect 6604 7352 6610 7404
rect 6638 7352 6644 7404
rect 6696 7352 6702 7404
rect 6914 7352 6920 7404
rect 6972 7352 6978 7404
rect 7006 7352 7012 7404
rect 7064 7392 7070 7404
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 7064 7364 7297 7392
rect 7064 7352 7070 7364
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 2608 7296 2774 7324
rect 1578 7148 1584 7200
rect 1636 7148 1642 7200
rect 2746 7188 2774 7296
rect 3234 7284 3240 7336
rect 3292 7324 3298 7336
rect 3694 7324 3700 7336
rect 3292 7296 3700 7324
rect 3292 7284 3298 7296
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 3789 7327 3847 7333
rect 3789 7293 3801 7327
rect 3835 7324 3847 7327
rect 4709 7327 4767 7333
rect 4709 7324 4721 7327
rect 3835 7296 4721 7324
rect 3835 7293 3847 7296
rect 3789 7287 3847 7293
rect 4709 7293 4721 7296
rect 4755 7293 4767 7327
rect 4709 7287 4767 7293
rect 4982 7284 4988 7336
rect 5040 7324 5046 7336
rect 5166 7324 5172 7336
rect 5040 7296 5172 7324
rect 5040 7284 5046 7296
rect 5166 7284 5172 7296
rect 5224 7324 5230 7336
rect 5445 7327 5503 7333
rect 5445 7324 5457 7327
rect 5224 7296 5457 7324
rect 5224 7284 5230 7296
rect 5445 7293 5457 7296
rect 5491 7293 5503 7327
rect 6380 7324 6408 7352
rect 7392 7324 7420 7355
rect 7466 7352 7472 7404
rect 7524 7352 7530 7404
rect 7668 7401 7696 7432
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 6380 7296 7420 7324
rect 5445 7287 5503 7293
rect 4617 7259 4675 7265
rect 4617 7225 4629 7259
rect 4663 7256 4675 7259
rect 5718 7256 5724 7268
rect 4663 7228 5724 7256
rect 4663 7225 4675 7228
rect 4617 7219 4675 7225
rect 5718 7216 5724 7228
rect 5776 7216 5782 7268
rect 3970 7188 3976 7200
rect 2746 7160 3976 7188
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 5902 7148 5908 7200
rect 5960 7188 5966 7200
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 5960 7160 6377 7188
rect 5960 7148 5966 7160
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 7098 7188 7104 7200
rect 6512 7160 7104 7188
rect 6512 7148 6518 7160
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 1104 7098 8096 7120
rect 1104 7046 1823 7098
rect 1875 7046 1887 7098
rect 1939 7046 1951 7098
rect 2003 7046 2015 7098
rect 2067 7046 2079 7098
rect 2131 7046 3570 7098
rect 3622 7046 3634 7098
rect 3686 7046 3698 7098
rect 3750 7046 3762 7098
rect 3814 7046 3826 7098
rect 3878 7046 5317 7098
rect 5369 7046 5381 7098
rect 5433 7046 5445 7098
rect 5497 7046 5509 7098
rect 5561 7046 5573 7098
rect 5625 7046 7064 7098
rect 7116 7046 7128 7098
rect 7180 7046 7192 7098
rect 7244 7046 7256 7098
rect 7308 7046 7320 7098
rect 7372 7046 8096 7098
rect 1104 7024 8096 7046
rect 1504 6956 1716 6984
rect 934 6808 940 6860
rect 992 6848 998 6860
rect 1504 6848 1532 6956
rect 1578 6876 1584 6928
rect 1636 6876 1642 6928
rect 1688 6925 1716 6956
rect 1762 6944 1768 6996
rect 1820 6984 1826 6996
rect 2314 6984 2320 6996
rect 1820 6956 2320 6984
rect 1820 6944 1826 6956
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 5629 6987 5687 6993
rect 5629 6953 5641 6987
rect 5675 6984 5687 6987
rect 5810 6984 5816 6996
rect 5675 6956 5816 6984
rect 5675 6953 5687 6956
rect 5629 6947 5687 6953
rect 5810 6944 5816 6956
rect 5868 6984 5874 6996
rect 5868 6956 7512 6984
rect 5868 6944 5874 6956
rect 1673 6919 1731 6925
rect 1673 6885 1685 6919
rect 1719 6885 1731 6919
rect 3142 6916 3148 6928
rect 1673 6879 1731 6885
rect 2608 6888 3148 6916
rect 992 6820 1532 6848
rect 992 6808 998 6820
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6780 1547 6783
rect 1596 6780 1624 6876
rect 1535 6752 1624 6780
rect 1535 6749 1547 6752
rect 1489 6743 1547 6749
rect 2406 6740 2412 6792
rect 2464 6740 2470 6792
rect 2498 6740 2504 6792
rect 2556 6789 2562 6792
rect 2556 6783 2579 6789
rect 2567 6780 2579 6783
rect 2608 6780 2636 6888
rect 3142 6876 3148 6888
rect 3200 6916 3206 6928
rect 3200 6888 4246 6916
rect 3200 6876 3206 6888
rect 2682 6808 2688 6860
rect 2740 6808 2746 6860
rect 3237 6851 3295 6857
rect 3237 6817 3249 6851
rect 3283 6848 3295 6851
rect 3418 6848 3424 6860
rect 3283 6820 3424 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 3510 6808 3516 6860
rect 3568 6848 3574 6860
rect 4218 6848 4246 6888
rect 7484 6860 7512 6956
rect 5350 6848 5356 6860
rect 3568 6820 4016 6848
rect 4218 6820 5356 6848
rect 3568 6808 3574 6820
rect 2567 6752 2636 6780
rect 2700 6780 2728 6808
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2700 6752 2789 6780
rect 2567 6749 2579 6752
rect 2556 6743 2579 6749
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6780 2927 6783
rect 2958 6780 2964 6792
rect 2915 6752 2964 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 2556 6740 2562 6743
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 3988 6789 4016 6820
rect 4264 6789 4292 6820
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 6638 6848 6644 6860
rect 5828 6820 6644 6848
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 2317 6715 2375 6721
rect 2317 6712 2329 6715
rect 1596 6684 2329 6712
rect 1486 6604 1492 6656
rect 1544 6644 1550 6656
rect 1596 6644 1624 6684
rect 2317 6681 2329 6684
rect 2363 6681 2375 6715
rect 2424 6712 2452 6740
rect 2685 6715 2743 6721
rect 2685 6712 2697 6715
rect 2424 6684 2697 6712
rect 2317 6675 2375 6681
rect 2685 6681 2697 6684
rect 2731 6681 2743 6715
rect 2685 6675 2743 6681
rect 3513 6715 3571 6721
rect 3513 6681 3525 6715
rect 3559 6712 3571 6715
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 3559 6684 3801 6712
rect 3559 6681 3571 6684
rect 3513 6675 3571 6681
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 3988 6712 4016 6743
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 4948 6752 5457 6780
rect 4948 6740 4954 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5074 6712 5080 6724
rect 3988 6684 5080 6712
rect 3789 6675 3847 6681
rect 5074 6672 5080 6684
rect 5132 6712 5138 6724
rect 5828 6712 5856 6820
rect 6638 6808 6644 6820
rect 6696 6808 6702 6860
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 7377 6851 7435 6857
rect 7377 6848 7389 6851
rect 6788 6820 7389 6848
rect 6788 6808 6794 6820
rect 7377 6817 7389 6820
rect 7423 6817 7435 6851
rect 7377 6811 7435 6817
rect 7466 6808 7472 6860
rect 7524 6808 7530 6860
rect 5132 6684 5856 6712
rect 5132 6672 5138 6684
rect 1544 6616 1624 6644
rect 1544 6604 1550 6616
rect 2222 6604 2228 6656
rect 2280 6604 2286 6656
rect 3050 6604 3056 6656
rect 3108 6604 3114 6656
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 4157 6647 4215 6653
rect 4157 6644 4169 6647
rect 4028 6616 4169 6644
rect 4028 6604 4034 6616
rect 4157 6613 4169 6616
rect 4203 6644 4215 6647
rect 4982 6644 4988 6656
rect 4203 6616 4988 6644
rect 4203 6613 4215 6616
rect 4157 6607 4215 6613
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5626 6644 5632 6656
rect 5307 6616 5632 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 6012 6644 6040 6766
rect 7101 6715 7159 6721
rect 7101 6681 7113 6715
rect 7147 6712 7159 6715
rect 7190 6712 7196 6724
rect 7147 6684 7196 6712
rect 7147 6681 7159 6684
rect 7101 6675 7159 6681
rect 7190 6672 7196 6684
rect 7248 6672 7254 6724
rect 5868 6616 6040 6644
rect 5868 6604 5874 6616
rect 1104 6554 8096 6576
rect 1104 6502 2483 6554
rect 2535 6502 2547 6554
rect 2599 6502 2611 6554
rect 2663 6502 2675 6554
rect 2727 6502 2739 6554
rect 2791 6502 4230 6554
rect 4282 6502 4294 6554
rect 4346 6502 4358 6554
rect 4410 6502 4422 6554
rect 4474 6502 4486 6554
rect 4538 6502 5977 6554
rect 6029 6502 6041 6554
rect 6093 6502 6105 6554
rect 6157 6502 6169 6554
rect 6221 6502 6233 6554
rect 6285 6502 7724 6554
rect 7776 6502 7788 6554
rect 7840 6502 7852 6554
rect 7904 6502 7916 6554
rect 7968 6502 7980 6554
rect 8032 6502 8096 6554
rect 1104 6480 8096 6502
rect 1394 6400 1400 6452
rect 1452 6400 1458 6452
rect 2866 6440 2872 6452
rect 1596 6412 2872 6440
rect 1596 6313 1624 6412
rect 2866 6400 2872 6412
rect 2924 6440 2930 6452
rect 3510 6440 3516 6452
rect 2924 6412 3516 6440
rect 2924 6400 2930 6412
rect 3510 6400 3516 6412
rect 3568 6400 3574 6452
rect 3651 6443 3709 6449
rect 3651 6409 3663 6443
rect 3697 6440 3709 6443
rect 3970 6440 3976 6452
rect 3697 6412 3976 6440
rect 3697 6409 3709 6412
rect 3651 6403 3709 6409
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 6472 6412 7512 6440
rect 3234 6332 3240 6384
rect 3292 6332 3298 6384
rect 4062 6372 4068 6384
rect 3804 6344 4068 6372
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1320 6276 1593 6304
rect 1320 6180 1348 6276
rect 1581 6273 1593 6276
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 1670 6264 1676 6316
rect 1728 6264 1734 6316
rect 1872 6276 2360 6304
rect 1872 6245 1900 6276
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6205 1915 6239
rect 1857 6199 1915 6205
rect 2222 6196 2228 6248
rect 2280 6196 2286 6248
rect 2332 6236 2360 6276
rect 2774 6236 2780 6248
rect 2332 6208 2780 6236
rect 2774 6196 2780 6208
rect 2832 6236 2838 6248
rect 3804 6245 3832 6344
rect 4062 6332 4068 6344
rect 4120 6332 4126 6384
rect 4706 6332 4712 6384
rect 4764 6332 4770 6384
rect 5368 6344 6408 6372
rect 5368 6316 5396 6344
rect 6380 6316 6408 6344
rect 6472 6316 6500 6412
rect 6549 6375 6607 6381
rect 6549 6341 6561 6375
rect 6595 6372 6607 6375
rect 7098 6372 7104 6384
rect 6595 6344 7104 6372
rect 6595 6341 6607 6344
rect 6549 6335 6607 6341
rect 7098 6332 7104 6344
rect 7156 6332 7162 6384
rect 7374 6332 7380 6384
rect 7432 6332 7438 6384
rect 5350 6264 5356 6316
rect 5408 6264 5414 6316
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 3789 6239 3847 6245
rect 3789 6236 3801 6239
rect 2832 6208 3801 6236
rect 2832 6196 2838 6208
rect 3789 6205 3801 6208
rect 3835 6205 3847 6239
rect 3789 6199 3847 6205
rect 4062 6196 4068 6248
rect 4120 6196 4126 6248
rect 4614 6196 4620 6248
rect 4672 6236 4678 6248
rect 5828 6236 5856 6267
rect 6362 6264 6368 6316
rect 6420 6264 6426 6316
rect 6454 6264 6460 6316
rect 6512 6304 6518 6316
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 6512 6276 6653 6304
rect 6512 6264 6518 6276
rect 6641 6273 6653 6276
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 4672 6208 5856 6236
rect 4672 6196 4678 6208
rect 1302 6128 1308 6180
rect 1360 6128 1366 6180
rect 3050 6128 3056 6180
rect 3108 6168 3114 6180
rect 3108 6140 3924 6168
rect 3108 6128 3114 6140
rect 2222 6060 2228 6112
rect 2280 6100 2286 6112
rect 3326 6100 3332 6112
rect 2280 6072 3332 6100
rect 2280 6060 2286 6072
rect 3326 6060 3332 6072
rect 3384 6060 3390 6112
rect 3896 6100 3924 6140
rect 6638 6128 6644 6180
rect 6696 6168 6702 6180
rect 6748 6168 6776 6267
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 6880 6276 7205 6304
rect 6880 6264 6886 6276
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6273 7343 6307
rect 7484 6304 7512 6412
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 7484 6276 7573 6304
rect 7285 6267 7343 6273
rect 7561 6273 7573 6276
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7300 6236 7328 6267
rect 8202 6236 8208 6248
rect 7156 6208 8208 6236
rect 7156 6196 7162 6208
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 6822 6168 6828 6180
rect 6696 6140 6828 6168
rect 6696 6128 6702 6140
rect 6822 6128 6828 6140
rect 6880 6128 6886 6180
rect 6917 6171 6975 6177
rect 6917 6137 6929 6171
rect 6963 6168 6975 6171
rect 7834 6168 7840 6180
rect 6963 6140 7840 6168
rect 6963 6137 6975 6140
rect 6917 6131 6975 6137
rect 7834 6128 7840 6140
rect 7892 6128 7898 6180
rect 5166 6100 5172 6112
rect 3896 6072 5172 6100
rect 5166 6060 5172 6072
rect 5224 6100 5230 6112
rect 5537 6103 5595 6109
rect 5537 6100 5549 6103
rect 5224 6072 5549 6100
rect 5224 6060 5230 6072
rect 5537 6069 5549 6072
rect 5583 6069 5595 6103
rect 5537 6063 5595 6069
rect 6089 6103 6147 6109
rect 6089 6069 6101 6103
rect 6135 6100 6147 6103
rect 6178 6100 6184 6112
rect 6135 6072 6184 6100
rect 6135 6069 6147 6072
rect 6089 6063 6147 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 7006 6060 7012 6112
rect 7064 6060 7070 6112
rect 7190 6060 7196 6112
rect 7248 6100 7254 6112
rect 7742 6100 7748 6112
rect 7248 6072 7748 6100
rect 7248 6060 7254 6072
rect 7742 6060 7748 6072
rect 7800 6060 7806 6112
rect 1104 6010 8096 6032
rect 1104 5958 1823 6010
rect 1875 5958 1887 6010
rect 1939 5958 1951 6010
rect 2003 5958 2015 6010
rect 2067 5958 2079 6010
rect 2131 5958 3570 6010
rect 3622 5958 3634 6010
rect 3686 5958 3698 6010
rect 3750 5958 3762 6010
rect 3814 5958 3826 6010
rect 3878 5958 5317 6010
rect 5369 5958 5381 6010
rect 5433 5958 5445 6010
rect 5497 5958 5509 6010
rect 5561 5958 5573 6010
rect 5625 5958 7064 6010
rect 7116 5958 7128 6010
rect 7180 5958 7192 6010
rect 7244 5958 7256 6010
rect 7308 5958 7320 6010
rect 7372 5958 8096 6010
rect 1104 5936 8096 5958
rect 1210 5856 1216 5908
rect 1268 5896 1274 5908
rect 1268 5868 3464 5896
rect 1268 5856 1274 5868
rect 1302 5788 1308 5840
rect 1360 5828 1366 5840
rect 2866 5828 2872 5840
rect 1360 5800 2872 5828
rect 1360 5788 1366 5800
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 1636 5732 2268 5760
rect 1636 5720 1642 5732
rect 1670 5652 1676 5704
rect 1728 5652 1734 5704
rect 2038 5652 2044 5704
rect 2096 5652 2102 5704
rect 2240 5701 2268 5732
rect 2424 5701 2452 5800
rect 2866 5788 2872 5800
rect 2924 5788 2930 5840
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 2648 5732 3280 5760
rect 2648 5720 2654 5732
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5661 2467 5695
rect 2409 5655 2467 5661
rect 2685 5671 2743 5677
rect 1302 5584 1308 5636
rect 1360 5624 1366 5636
rect 1688 5624 1716 5652
rect 2685 5637 2697 5671
rect 2731 5668 2743 5671
rect 2731 5640 2820 5668
rect 3050 5652 3056 5704
rect 3108 5652 3114 5704
rect 3142 5652 3148 5704
rect 3200 5652 3206 5704
rect 3252 5701 3280 5732
rect 3436 5701 3464 5868
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 4120 5868 4445 5896
rect 4120 5856 4126 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 4982 5856 4988 5908
rect 5040 5896 5046 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 5040 5868 5365 5896
rect 5040 5856 5046 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 6454 5896 6460 5908
rect 5353 5859 5411 5865
rect 5736 5868 6460 5896
rect 5736 5828 5764 5868
rect 6454 5856 6460 5868
rect 6512 5856 6518 5908
rect 7653 5899 7711 5905
rect 7653 5865 7665 5899
rect 7699 5896 7711 5899
rect 8110 5896 8116 5908
rect 7699 5868 8116 5896
rect 7699 5865 7711 5868
rect 7653 5859 7711 5865
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 3896 5800 5764 5828
rect 3896 5701 3924 5800
rect 7374 5788 7380 5840
rect 7432 5828 7438 5840
rect 7742 5828 7748 5840
rect 7432 5800 7748 5828
rect 7432 5788 7438 5800
rect 7742 5788 7748 5800
rect 7800 5788 7806 5840
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5760 5687 5763
rect 6638 5760 6644 5772
rect 5675 5732 6644 5760
rect 5675 5729 5687 5732
rect 5629 5723 5687 5729
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 3881 5695 3939 5701
rect 3881 5692 3893 5695
rect 3467 5664 3893 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 3881 5661 3893 5664
rect 3927 5661 3939 5695
rect 3881 5655 3939 5661
rect 3970 5652 3976 5704
rect 4028 5692 4034 5704
rect 4985 5695 5043 5701
rect 4985 5692 4997 5695
rect 4028 5664 4997 5692
rect 4028 5652 4034 5664
rect 4985 5661 4997 5664
rect 5031 5692 5043 5695
rect 5169 5695 5227 5701
rect 5169 5692 5181 5695
rect 5031 5664 5181 5692
rect 5031 5661 5043 5664
rect 4985 5655 5043 5661
rect 5169 5661 5181 5664
rect 5215 5661 5227 5695
rect 5169 5655 5227 5661
rect 7469 5695 7527 5701
rect 7469 5661 7481 5695
rect 7515 5692 7527 5695
rect 7834 5692 7840 5704
rect 7515 5664 7840 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 2731 5637 2743 5640
rect 2133 5627 2191 5633
rect 2685 5631 2743 5637
rect 2133 5624 2145 5627
rect 1360 5596 2145 5624
rect 1360 5584 1366 5596
rect 2133 5593 2145 5596
rect 2179 5593 2191 5627
rect 2792 5624 2820 5640
rect 2133 5587 2191 5593
rect 2240 5596 2636 5624
rect 2792 5596 3188 5624
rect 1670 5516 1676 5568
rect 1728 5556 1734 5568
rect 1857 5559 1915 5565
rect 1857 5556 1869 5559
rect 1728 5528 1869 5556
rect 1728 5516 1734 5528
rect 1857 5525 1869 5528
rect 1903 5525 1915 5559
rect 1857 5519 1915 5525
rect 2038 5516 2044 5568
rect 2096 5556 2102 5568
rect 2240 5556 2268 5596
rect 2096 5528 2268 5556
rect 2096 5516 2102 5528
rect 2406 5516 2412 5568
rect 2464 5556 2470 5568
rect 2501 5559 2559 5565
rect 2501 5556 2513 5559
rect 2464 5528 2513 5556
rect 2464 5516 2470 5528
rect 2501 5525 2513 5528
rect 2547 5525 2559 5559
rect 2608 5556 2636 5596
rect 2869 5559 2927 5565
rect 2869 5556 2881 5559
rect 2608 5528 2881 5556
rect 2501 5519 2559 5525
rect 2869 5525 2881 5528
rect 2915 5525 2927 5559
rect 3160 5556 3188 5596
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 4249 5627 4307 5633
rect 4249 5624 4261 5627
rect 4212 5596 4261 5624
rect 4212 5584 4218 5596
rect 4249 5593 4261 5596
rect 4295 5593 4307 5627
rect 4249 5587 4307 5593
rect 4706 5584 4712 5636
rect 4764 5584 4770 5636
rect 5902 5584 5908 5636
rect 5960 5584 5966 5636
rect 6012 5596 6394 5624
rect 3234 5556 3240 5568
rect 3160 5528 3240 5556
rect 2869 5519 2927 5525
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 4724 5556 4752 5584
rect 5166 5556 5172 5568
rect 4724 5528 5172 5556
rect 5166 5516 5172 5528
rect 5224 5556 5230 5568
rect 6012 5556 6040 5596
rect 5224 5528 6040 5556
rect 5224 5516 5230 5528
rect 6178 5516 6184 5568
rect 6236 5556 6242 5568
rect 6638 5556 6644 5568
rect 6236 5528 6644 5556
rect 6236 5516 6242 5528
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 6822 5516 6828 5568
rect 6880 5556 6886 5568
rect 7377 5559 7435 5565
rect 7377 5556 7389 5559
rect 6880 5528 7389 5556
rect 6880 5516 6886 5528
rect 7377 5525 7389 5528
rect 7423 5525 7435 5559
rect 7377 5519 7435 5525
rect 1104 5466 8096 5488
rect 1104 5414 2483 5466
rect 2535 5414 2547 5466
rect 2599 5414 2611 5466
rect 2663 5414 2675 5466
rect 2727 5414 2739 5466
rect 2791 5414 4230 5466
rect 4282 5414 4294 5466
rect 4346 5414 4358 5466
rect 4410 5414 4422 5466
rect 4474 5414 4486 5466
rect 4538 5414 5977 5466
rect 6029 5414 6041 5466
rect 6093 5414 6105 5466
rect 6157 5414 6169 5466
rect 6221 5414 6233 5466
rect 6285 5414 7724 5466
rect 7776 5414 7788 5466
rect 7840 5414 7852 5466
rect 7904 5414 7916 5466
rect 7968 5414 7980 5466
rect 8032 5414 8096 5466
rect 1104 5392 8096 5414
rect 2222 5312 2228 5364
rect 2280 5352 2286 5364
rect 2280 5324 2636 5352
rect 2280 5312 2286 5324
rect 1765 5287 1823 5293
rect 1765 5253 1777 5287
rect 1811 5284 1823 5287
rect 2038 5284 2044 5296
rect 1811 5256 2044 5284
rect 1811 5253 1823 5256
rect 1765 5247 1823 5253
rect 2038 5244 2044 5256
rect 2096 5244 2102 5296
rect 2608 5293 2636 5324
rect 3970 5312 3976 5364
rect 4028 5312 4034 5364
rect 6362 5312 6368 5364
rect 6420 5352 6426 5364
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 6420 5324 6469 5352
rect 6420 5312 6426 5324
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 6825 5355 6883 5361
rect 6825 5321 6837 5355
rect 6871 5352 6883 5355
rect 7466 5352 7472 5364
rect 6871 5324 7472 5352
rect 6871 5321 6883 5324
rect 6825 5315 6883 5321
rect 7466 5312 7472 5324
rect 7524 5312 7530 5364
rect 2593 5287 2651 5293
rect 2593 5253 2605 5287
rect 2639 5253 2651 5287
rect 2593 5247 2651 5253
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 1949 5219 2007 5225
rect 1949 5216 1961 5219
rect 1636 5188 1961 5216
rect 1636 5176 1642 5188
rect 1949 5185 1961 5188
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2385 5219 2443 5225
rect 2385 5185 2397 5219
rect 2431 5216 2443 5219
rect 2431 5185 2452 5216
rect 2385 5179 2452 5185
rect 1302 5108 1308 5160
rect 1360 5108 1366 5160
rect 2424 5148 2452 5179
rect 2498 5176 2504 5228
rect 2556 5176 2562 5228
rect 2774 5176 2780 5228
rect 2832 5176 2838 5228
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5216 3019 5219
rect 3326 5216 3332 5228
rect 3007 5188 3332 5216
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5185 3939 5219
rect 3988 5216 4016 5312
rect 6181 5287 6239 5293
rect 6181 5253 6193 5287
rect 6227 5284 6239 5287
rect 7650 5284 7656 5296
rect 6227 5256 7656 5284
rect 6227 5253 6239 5256
rect 6181 5247 6239 5253
rect 7650 5244 7656 5256
rect 7708 5244 7714 5296
rect 6641 5219 6699 5225
rect 3988 5188 4108 5216
rect 3881 5179 3939 5185
rect 3050 5148 3056 5160
rect 2424 5120 3056 5148
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 1320 5080 1348 5108
rect 2498 5080 2504 5092
rect 1320 5052 2504 5080
rect 2498 5040 2504 5052
rect 2556 5040 2562 5092
rect 3142 5040 3148 5092
rect 3200 5040 3206 5092
rect 934 4972 940 5024
rect 992 5012 998 5024
rect 1489 5015 1547 5021
rect 1489 5012 1501 5015
rect 992 4984 1501 5012
rect 992 4972 998 4984
rect 1489 4981 1501 4984
rect 1535 4981 1547 5015
rect 1489 4975 1547 4981
rect 2130 4972 2136 5024
rect 2188 4972 2194 5024
rect 2222 4972 2228 5024
rect 2280 4972 2286 5024
rect 3050 4972 3056 5024
rect 3108 5012 3114 5024
rect 3513 5015 3571 5021
rect 3513 5012 3525 5015
rect 3108 4984 3525 5012
rect 3108 4972 3114 4984
rect 3513 4981 3525 4984
rect 3559 4981 3571 5015
rect 3896 5012 3924 5179
rect 4080 5157 4108 5188
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 3973 5151 4031 5157
rect 3973 5117 3985 5151
rect 4019 5117 4031 5151
rect 3973 5111 4031 5117
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5117 4123 5151
rect 4065 5111 4123 5117
rect 3988 5080 4016 5111
rect 5902 5080 5908 5092
rect 3988 5052 5908 5080
rect 5902 5040 5908 5052
rect 5960 5080 5966 5092
rect 6656 5080 6684 5179
rect 7374 5176 7380 5228
rect 7432 5176 7438 5228
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5216 7803 5219
rect 8110 5216 8116 5228
rect 7791 5188 8116 5216
rect 7791 5185 7803 5188
rect 7745 5179 7803 5185
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 5960 5052 6684 5080
rect 5960 5040 5966 5052
rect 4154 5012 4160 5024
rect 3896 4984 4160 5012
rect 3513 4975 3571 4981
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 4709 5015 4767 5021
rect 4709 5012 4721 5015
rect 4672 4984 4721 5012
rect 4672 4972 4678 4984
rect 4709 4981 4721 4984
rect 4755 4981 4767 5015
rect 4709 4975 4767 4981
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 7561 5015 7619 5021
rect 7561 5012 7573 5015
rect 5868 4984 7573 5012
rect 5868 4972 5874 4984
rect 7561 4981 7573 4984
rect 7607 5012 7619 5015
rect 7650 5012 7656 5024
rect 7607 4984 7656 5012
rect 7607 4981 7619 4984
rect 7561 4975 7619 4981
rect 7650 4972 7656 4984
rect 7708 4972 7714 5024
rect 1104 4922 8096 4944
rect 1104 4870 1823 4922
rect 1875 4870 1887 4922
rect 1939 4870 1951 4922
rect 2003 4870 2015 4922
rect 2067 4870 2079 4922
rect 2131 4870 3570 4922
rect 3622 4870 3634 4922
rect 3686 4870 3698 4922
rect 3750 4870 3762 4922
rect 3814 4870 3826 4922
rect 3878 4870 5317 4922
rect 5369 4870 5381 4922
rect 5433 4870 5445 4922
rect 5497 4870 5509 4922
rect 5561 4870 5573 4922
rect 5625 4870 7064 4922
rect 7116 4870 7128 4922
rect 7180 4870 7192 4922
rect 7244 4870 7256 4922
rect 7308 4870 7320 4922
rect 7372 4870 8096 4922
rect 1104 4848 8096 4870
rect 3050 4768 3056 4820
rect 3108 4768 3114 4820
rect 4525 4811 4583 4817
rect 4525 4777 4537 4811
rect 4571 4808 4583 4811
rect 4890 4808 4896 4820
rect 4571 4780 4896 4808
rect 4571 4777 4583 4780
rect 4525 4771 4583 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 6730 4768 6736 4820
rect 6788 4768 6794 4820
rect 2593 4743 2651 4749
rect 2593 4709 2605 4743
rect 2639 4740 2651 4743
rect 2866 4740 2872 4752
rect 2639 4712 2872 4740
rect 2639 4709 2651 4712
rect 2593 4703 2651 4709
rect 2866 4700 2872 4712
rect 2924 4700 2930 4752
rect 3068 4740 3096 4768
rect 4154 4740 4160 4752
rect 2976 4712 3096 4740
rect 3896 4712 4160 4740
rect 2222 4632 2228 4684
rect 2280 4632 2286 4684
rect 1670 4564 1676 4616
rect 1728 4604 1734 4616
rect 1765 4607 1823 4613
rect 1765 4604 1777 4607
rect 1728 4576 1777 4604
rect 1728 4564 1734 4576
rect 1765 4573 1777 4576
rect 1811 4573 1823 4607
rect 2240 4604 2268 4632
rect 2317 4607 2375 4613
rect 2317 4604 2329 4607
rect 2240 4576 2329 4604
rect 1765 4567 1823 4573
rect 2317 4573 2329 4576
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4604 2835 4607
rect 2976 4604 3004 4712
rect 3421 4675 3479 4681
rect 3421 4672 3433 4675
rect 2823 4576 3004 4604
rect 3068 4644 3433 4672
rect 2823 4573 2835 4576
rect 2777 4567 2835 4573
rect 1394 4496 1400 4548
rect 1452 4496 1458 4548
rect 1946 4496 1952 4548
rect 2004 4496 2010 4548
rect 2038 4496 2044 4548
rect 2096 4536 2102 4548
rect 3068 4536 3096 4644
rect 3421 4641 3433 4644
rect 3467 4641 3479 4675
rect 3421 4635 3479 4641
rect 3234 4564 3240 4616
rect 3292 4564 3298 4616
rect 3252 4536 3280 4564
rect 2096 4508 3096 4536
rect 3160 4508 3280 4536
rect 2096 4496 2102 4508
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 3160 4468 3188 4508
rect 3896 4480 3924 4712
rect 4154 4700 4160 4712
rect 4212 4700 4218 4752
rect 3970 4632 3976 4684
rect 4028 4632 4034 4684
rect 6362 4672 6368 4684
rect 4172 4644 6368 4672
rect 4172 4613 4200 4644
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 7466 4672 7472 4684
rect 6880 4644 7472 4672
rect 6880 4632 6886 4644
rect 7466 4632 7472 4644
rect 7524 4672 7530 4684
rect 7653 4675 7711 4681
rect 7653 4672 7665 4675
rect 7524 4644 7665 4672
rect 7524 4632 7530 4644
rect 7653 4641 7665 4644
rect 7699 4641 7711 4675
rect 7653 4635 7711 4641
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4573 4215 4607
rect 4157 4567 4215 4573
rect 4522 4564 4528 4616
rect 4580 4564 4586 4616
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 4632 4576 5273 4604
rect 4065 4539 4123 4545
rect 4065 4505 4077 4539
rect 4111 4536 4123 4539
rect 4540 4536 4568 4564
rect 4632 4548 4660 4576
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 4111 4508 4568 4536
rect 4111 4505 4123 4508
rect 4065 4499 4123 4505
rect 4614 4496 4620 4548
rect 4672 4496 4678 4548
rect 4801 4539 4859 4545
rect 4801 4505 4813 4539
rect 4847 4505 4859 4539
rect 4801 4499 4859 4505
rect 5169 4539 5227 4545
rect 5169 4505 5181 4539
rect 5215 4536 5227 4539
rect 8386 4536 8392 4548
rect 5215 4508 8392 4536
rect 5215 4505 5227 4508
rect 5169 4499 5227 4505
rect 2915 4440 3188 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 3234 4428 3240 4480
rect 3292 4428 3298 4480
rect 3329 4471 3387 4477
rect 3329 4437 3341 4471
rect 3375 4468 3387 4471
rect 3878 4468 3884 4480
rect 3375 4440 3884 4468
rect 3375 4437 3387 4440
rect 3329 4431 3387 4437
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4816 4468 4844 4499
rect 8386 4496 8392 4508
rect 8444 4496 8450 4548
rect 4212 4440 4844 4468
rect 4212 4428 4218 4440
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 7101 4471 7159 4477
rect 7101 4468 7113 4471
rect 5868 4440 7113 4468
rect 5868 4428 5874 4440
rect 7101 4437 7113 4440
rect 7147 4437 7159 4471
rect 7101 4431 7159 4437
rect 1104 4378 8096 4400
rect 1104 4326 2483 4378
rect 2535 4326 2547 4378
rect 2599 4326 2611 4378
rect 2663 4326 2675 4378
rect 2727 4326 2739 4378
rect 2791 4326 4230 4378
rect 4282 4326 4294 4378
rect 4346 4326 4358 4378
rect 4410 4326 4422 4378
rect 4474 4326 4486 4378
rect 4538 4326 5977 4378
rect 6029 4326 6041 4378
rect 6093 4326 6105 4378
rect 6157 4326 6169 4378
rect 6221 4326 6233 4378
rect 6285 4326 7724 4378
rect 7776 4326 7788 4378
rect 7840 4326 7852 4378
rect 7904 4326 7916 4378
rect 7968 4326 7980 4378
rect 8032 4326 8096 4378
rect 1104 4304 8096 4326
rect 1302 4224 1308 4276
rect 1360 4224 1366 4276
rect 1578 4224 1584 4276
rect 1636 4264 1642 4276
rect 3418 4264 3424 4276
rect 1636 4236 3424 4264
rect 1636 4224 1642 4236
rect 3418 4224 3424 4236
rect 3476 4224 3482 4276
rect 5626 4264 5632 4276
rect 4632 4236 5632 4264
rect 1320 4196 1348 4224
rect 4246 4196 4252 4208
rect 1320 4168 2176 4196
rect 3818 4168 4252 4196
rect 1210 4088 1216 4140
rect 1268 4128 1274 4140
rect 1857 4131 1915 4137
rect 1857 4128 1869 4131
rect 1268 4100 1869 4128
rect 1268 4088 1274 4100
rect 1596 4072 1624 4100
rect 1857 4097 1869 4100
rect 1903 4097 1915 4131
rect 1857 4091 1915 4097
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4128 2007 4131
rect 2038 4128 2044 4140
rect 1995 4100 2044 4128
rect 1995 4097 2007 4100
rect 1949 4091 2007 4097
rect 1578 4020 1584 4072
rect 1636 4020 1642 4072
rect 1670 4020 1676 4072
rect 1728 4060 1734 4072
rect 1964 4060 1992 4091
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 2148 4137 2176 4168
rect 4246 4156 4252 4168
rect 4304 4156 4310 4208
rect 4632 4205 4660 4236
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 5902 4224 5908 4276
rect 5960 4264 5966 4276
rect 6089 4267 6147 4273
rect 6089 4264 6101 4267
rect 5960 4236 6101 4264
rect 5960 4224 5966 4236
rect 6089 4233 6101 4236
rect 6135 4233 6147 4267
rect 6089 4227 6147 4233
rect 4617 4199 4675 4205
rect 4617 4165 4629 4199
rect 4663 4165 4675 4199
rect 4617 4159 4675 4165
rect 5166 4156 5172 4208
rect 5224 4156 5230 4208
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4097 2191 4131
rect 4341 4131 4399 4137
rect 2133 4091 2191 4097
rect 2424 4100 2912 4128
rect 1728 4032 1992 4060
rect 1728 4020 1734 4032
rect 2222 4020 2228 4072
rect 2280 4060 2286 4072
rect 2424 4069 2452 4100
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 2280 4032 2421 4060
rect 2280 4020 2286 4032
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 2774 4020 2780 4072
rect 2832 4020 2838 4072
rect 2884 4060 2912 4100
rect 4341 4097 4353 4131
rect 4387 4097 4399 4131
rect 6104 4128 6132 4227
rect 6362 4224 6368 4276
rect 6420 4224 6426 4276
rect 7466 4224 7472 4276
rect 7524 4224 7530 4276
rect 7558 4224 7564 4276
rect 7616 4264 7622 4276
rect 7745 4267 7803 4273
rect 7745 4264 7757 4267
rect 7616 4236 7757 4264
rect 7616 4224 7622 4236
rect 7745 4233 7757 4236
rect 7791 4233 7803 4267
rect 7745 4227 7803 4233
rect 7374 4156 7380 4208
rect 7432 4156 7438 4208
rect 7484 4196 7512 4224
rect 7484 4168 7604 4196
rect 7576 4137 7604 4168
rect 8202 4156 8208 4208
rect 8260 4156 8266 4208
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 6104 4100 6929 4128
rect 4341 4091 4399 4097
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4128 7619 4131
rect 7742 4128 7748 4140
rect 7607 4100 7748 4128
rect 7607 4097 7619 4100
rect 7561 4091 7619 4097
rect 2958 4060 2964 4072
rect 2884 4032 2964 4060
rect 2958 4020 2964 4032
rect 3016 4060 3022 4072
rect 4356 4060 4384 4091
rect 3016 4032 4384 4060
rect 3016 4020 3022 4032
rect 6454 4020 6460 4072
rect 6512 4060 6518 4072
rect 6822 4060 6828 4072
rect 6512 4032 6828 4060
rect 6512 4020 6518 4032
rect 6822 4020 6828 4032
rect 6880 4060 6886 4072
rect 7208 4060 7236 4091
rect 6880 4032 7236 4060
rect 7484 4060 7512 4091
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 7834 4060 7840 4072
rect 7484 4032 7840 4060
rect 6880 4020 6886 4032
rect 7834 4020 7840 4032
rect 7892 4060 7898 4072
rect 8220 4060 8248 4156
rect 7892 4032 8248 4060
rect 7892 4020 7898 4032
rect 14 3884 20 3936
rect 72 3924 78 3936
rect 1946 3924 1952 3936
rect 72 3896 1952 3924
rect 72 3884 78 3896
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 3326 3924 3332 3936
rect 2363 3896 3332 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 3326 3884 3332 3896
rect 3384 3884 3390 3936
rect 3878 3884 3884 3936
rect 3936 3924 3942 3936
rect 4203 3927 4261 3933
rect 4203 3924 4215 3927
rect 3936 3896 4215 3924
rect 3936 3884 3942 3896
rect 4203 3893 4215 3896
rect 4249 3924 4261 3927
rect 5074 3924 5080 3936
rect 4249 3896 5080 3924
rect 4249 3893 4261 3896
rect 4203 3887 4261 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 7650 3924 7656 3936
rect 6512 3896 7656 3924
rect 6512 3884 6518 3896
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 1104 3834 8096 3856
rect 1104 3782 1823 3834
rect 1875 3782 1887 3834
rect 1939 3782 1951 3834
rect 2003 3782 2015 3834
rect 2067 3782 2079 3834
rect 2131 3782 3570 3834
rect 3622 3782 3634 3834
rect 3686 3782 3698 3834
rect 3750 3782 3762 3834
rect 3814 3782 3826 3834
rect 3878 3782 5317 3834
rect 5369 3782 5381 3834
rect 5433 3782 5445 3834
rect 5497 3782 5509 3834
rect 5561 3782 5573 3834
rect 5625 3782 7064 3834
rect 7116 3782 7128 3834
rect 7180 3782 7192 3834
rect 7244 3782 7256 3834
rect 7308 3782 7320 3834
rect 7372 3782 8096 3834
rect 1104 3760 8096 3782
rect 1486 3680 1492 3732
rect 1544 3720 1550 3732
rect 6362 3720 6368 3732
rect 1544 3692 6368 3720
rect 1544 3680 1550 3692
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 7558 3680 7564 3732
rect 7616 3720 7622 3732
rect 7653 3723 7711 3729
rect 7653 3720 7665 3723
rect 7616 3692 7665 3720
rect 7616 3680 7622 3692
rect 7653 3689 7665 3692
rect 7699 3689 7711 3723
rect 7653 3683 7711 3689
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 2222 3584 2228 3596
rect 1903 3556 2228 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 4246 3584 4252 3596
rect 2924 3556 4252 3584
rect 2924 3544 2930 3556
rect 3252 3502 3280 3556
rect 4246 3544 4252 3556
rect 4304 3584 4310 3596
rect 5166 3584 5172 3596
rect 4304 3556 5172 3584
rect 4304 3544 4310 3556
rect 3786 3476 3792 3528
rect 3844 3476 3850 3528
rect 4062 3476 4068 3528
rect 4120 3476 4126 3528
rect 4448 3502 4476 3556
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 5813 3587 5871 3593
rect 5813 3553 5825 3587
rect 5859 3584 5871 3587
rect 5905 3587 5963 3593
rect 5905 3584 5917 3587
rect 5859 3556 5917 3584
rect 5859 3553 5871 3556
rect 5813 3547 5871 3553
rect 5905 3553 5917 3556
rect 5951 3584 5963 3587
rect 6730 3584 6736 3596
rect 5951 3556 6736 3584
rect 5951 3553 5963 3556
rect 5905 3547 5963 3553
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 2133 3451 2191 3457
rect 2133 3417 2145 3451
rect 2179 3448 2191 3451
rect 2406 3448 2412 3460
rect 2179 3420 2412 3448
rect 2179 3417 2191 3420
rect 2133 3411 2191 3417
rect 2406 3408 2412 3420
rect 2464 3408 2470 3460
rect 4080 3448 4108 3476
rect 3620 3420 4108 3448
rect 5537 3451 5595 3457
rect 3620 3392 3648 3420
rect 5537 3417 5549 3451
rect 5583 3448 5595 3451
rect 5810 3448 5816 3460
rect 5583 3420 5816 3448
rect 5583 3417 5595 3420
rect 5537 3411 5595 3417
rect 5810 3408 5816 3420
rect 5868 3408 5874 3460
rect 5902 3408 5908 3460
rect 5960 3448 5966 3460
rect 6181 3451 6239 3457
rect 6181 3448 6193 3451
rect 5960 3420 6193 3448
rect 5960 3408 5966 3420
rect 6181 3417 6193 3420
rect 6227 3417 6239 3451
rect 6181 3411 6239 3417
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 6512 3420 6670 3448
rect 6512 3408 6518 3420
rect 7466 3408 7472 3460
rect 7524 3448 7530 3460
rect 7742 3448 7748 3460
rect 7524 3420 7748 3448
rect 7524 3408 7530 3420
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 7834 3408 7840 3460
rect 7892 3408 7898 3460
rect 3142 3340 3148 3392
rect 3200 3380 3206 3392
rect 3602 3380 3608 3392
rect 3200 3352 3608 3380
rect 3200 3340 3206 3352
rect 3602 3340 3608 3352
rect 3660 3340 3666 3392
rect 3970 3340 3976 3392
rect 4028 3340 4034 3392
rect 4065 3383 4123 3389
rect 4065 3349 4077 3383
rect 4111 3380 4123 3383
rect 5258 3380 5264 3392
rect 4111 3352 5264 3380
rect 4111 3349 4123 3352
rect 4065 3343 4123 3349
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 7098 3340 7104 3392
rect 7156 3380 7162 3392
rect 7852 3380 7880 3408
rect 7156 3352 7880 3380
rect 7156 3340 7162 3352
rect 1104 3290 8096 3312
rect 1104 3238 2483 3290
rect 2535 3238 2547 3290
rect 2599 3238 2611 3290
rect 2663 3238 2675 3290
rect 2727 3238 2739 3290
rect 2791 3238 4230 3290
rect 4282 3238 4294 3290
rect 4346 3238 4358 3290
rect 4410 3238 4422 3290
rect 4474 3238 4486 3290
rect 4538 3238 5977 3290
rect 6029 3238 6041 3290
rect 6093 3238 6105 3290
rect 6157 3238 6169 3290
rect 6221 3238 6233 3290
rect 6285 3238 7724 3290
rect 7776 3238 7788 3290
rect 7840 3238 7852 3290
rect 7904 3238 7916 3290
rect 7968 3238 7980 3290
rect 8032 3238 8096 3290
rect 1104 3216 8096 3238
rect 1670 3136 1676 3188
rect 1728 3176 1734 3188
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 1728 3148 2145 3176
rect 1728 3136 1734 3148
rect 2133 3145 2145 3148
rect 2179 3176 2191 3179
rect 2406 3176 2412 3188
rect 2179 3148 2412 3176
rect 2179 3145 2191 3148
rect 2133 3139 2191 3145
rect 2406 3136 2412 3148
rect 2464 3136 2470 3188
rect 2501 3179 2559 3185
rect 2501 3145 2513 3179
rect 2547 3176 2559 3179
rect 2547 3148 3372 3176
rect 2547 3145 2559 3148
rect 2501 3139 2559 3145
rect 3344 3108 3372 3148
rect 3418 3136 3424 3188
rect 3476 3176 3482 3188
rect 4433 3179 4491 3185
rect 4433 3176 4445 3179
rect 3476 3148 4445 3176
rect 3476 3136 3482 3148
rect 4433 3145 4445 3148
rect 4479 3145 4491 3179
rect 4433 3139 4491 3145
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 4801 3179 4859 3185
rect 4801 3176 4813 3179
rect 4764 3148 4813 3176
rect 4764 3136 4770 3148
rect 4801 3145 4813 3148
rect 4847 3145 4859 3179
rect 4801 3139 4859 3145
rect 5902 3136 5908 3188
rect 5960 3136 5966 3188
rect 6362 3136 6368 3188
rect 6420 3176 6426 3188
rect 7101 3179 7159 3185
rect 7101 3176 7113 3179
rect 6420 3148 7113 3176
rect 6420 3136 6426 3148
rect 7101 3145 7113 3148
rect 7147 3145 7159 3179
rect 7101 3139 7159 3145
rect 7466 3136 7472 3188
rect 7524 3136 7530 3188
rect 4154 3108 4160 3120
rect 1872 3080 2728 3108
rect 3344 3080 4160 3108
rect 1872 3049 1900 3080
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2038 3000 2044 3052
rect 2096 3000 2102 3052
rect 2317 3043 2375 3049
rect 2317 3040 2329 3043
rect 2148 3012 2329 3040
rect 1578 2932 1584 2984
rect 1636 2972 1642 2984
rect 2148 2972 2176 3012
rect 2317 3009 2329 3012
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 1636 2944 2176 2972
rect 1636 2932 1642 2944
rect 2222 2932 2228 2984
rect 2280 2972 2286 2984
rect 2593 2975 2651 2981
rect 2593 2972 2605 2975
rect 2280 2944 2605 2972
rect 2280 2932 2286 2944
rect 2593 2941 2605 2944
rect 2639 2941 2651 2975
rect 2700 2972 2728 3080
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 4614 3108 4620 3120
rect 4387 3080 4620 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 4614 3068 4620 3080
rect 4672 3068 4678 3120
rect 6546 3068 6552 3120
rect 6604 3068 6610 3120
rect 6822 3068 6828 3120
rect 6880 3108 6886 3120
rect 7484 3108 7512 3136
rect 6880 3080 7236 3108
rect 6880 3068 6886 3080
rect 5258 3000 5264 3052
rect 5316 3040 5322 3052
rect 5718 3040 5724 3052
rect 5316 3012 5724 3040
rect 5316 3000 5322 3012
rect 5718 3000 5724 3012
rect 5776 3040 5782 3052
rect 6733 3043 6791 3049
rect 6733 3040 6745 3043
rect 5776 3012 6745 3040
rect 5776 3000 5782 3012
rect 6733 3009 6745 3012
rect 6779 3009 6791 3043
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 6733 3003 6791 3009
rect 6840 3012 7021 3040
rect 3418 2972 3424 2984
rect 2700 2944 3424 2972
rect 2593 2935 2651 2941
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 3602 2932 3608 2984
rect 3660 2972 3666 2984
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 3660 2944 4905 2972
rect 3660 2932 3666 2944
rect 4893 2941 4905 2944
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 4982 2932 4988 2984
rect 5040 2932 5046 2984
rect 5166 2932 5172 2984
rect 5224 2972 5230 2984
rect 6840 2972 6868 3012
rect 7009 3009 7021 3012
rect 7055 3040 7067 3043
rect 7098 3040 7104 3052
rect 7055 3012 7104 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 5224 2944 6868 2972
rect 6917 2975 6975 2981
rect 5224 2932 5230 2944
rect 6917 2941 6929 2975
rect 6963 2972 6975 2975
rect 7208 2972 7236 3080
rect 7300 3080 7512 3108
rect 7300 3049 7328 3080
rect 7558 3068 7564 3120
rect 7616 3068 7622 3120
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3040 7527 3043
rect 7576 3040 7604 3068
rect 7515 3012 7604 3040
rect 7515 3009 7527 3012
rect 7469 3003 7527 3009
rect 6963 2944 7236 2972
rect 6963 2941 6975 2944
rect 6917 2935 6975 2941
rect 1780 2876 2636 2904
rect 1780 2845 1808 2876
rect 1765 2839 1823 2845
rect 1765 2805 1777 2839
rect 1811 2805 1823 2839
rect 2608 2836 2636 2876
rect 2682 2864 2688 2916
rect 2740 2904 2746 2916
rect 4246 2904 4252 2916
rect 2740 2876 4252 2904
rect 2740 2864 2746 2876
rect 4246 2864 4252 2876
rect 4304 2904 4310 2916
rect 5000 2904 5028 2932
rect 4304 2876 5028 2904
rect 4304 2864 4310 2876
rect 4154 2836 4160 2848
rect 2608 2808 4160 2836
rect 1765 2799 1823 2805
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 6822 2796 6828 2848
rect 6880 2836 6886 2848
rect 7392 2836 7420 3003
rect 7650 3000 7656 3052
rect 7708 3000 7714 3052
rect 6880 2808 7420 2836
rect 6880 2796 6886 2808
rect 1104 2746 8096 2768
rect 1104 2694 1823 2746
rect 1875 2694 1887 2746
rect 1939 2694 1951 2746
rect 2003 2694 2015 2746
rect 2067 2694 2079 2746
rect 2131 2694 3570 2746
rect 3622 2694 3634 2746
rect 3686 2694 3698 2746
rect 3750 2694 3762 2746
rect 3814 2694 3826 2746
rect 3878 2694 5317 2746
rect 5369 2694 5381 2746
rect 5433 2694 5445 2746
rect 5497 2694 5509 2746
rect 5561 2694 5573 2746
rect 5625 2694 7064 2746
rect 7116 2694 7128 2746
rect 7180 2694 7192 2746
rect 7244 2694 7256 2746
rect 7308 2694 7320 2746
rect 7372 2694 8096 2746
rect 1104 2672 8096 2694
rect 3789 2635 3847 2641
rect 3789 2601 3801 2635
rect 3835 2632 3847 2635
rect 3970 2632 3976 2644
rect 3835 2604 3976 2632
rect 3835 2601 3847 2604
rect 3789 2595 3847 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 5166 2592 5172 2644
rect 5224 2592 5230 2644
rect 5718 2592 5724 2644
rect 5776 2592 5782 2644
rect 7650 2592 7656 2644
rect 7708 2592 7714 2644
rect 3605 2567 3663 2573
rect 3605 2533 3617 2567
rect 3651 2533 3663 2567
rect 5184 2564 5212 2592
rect 5736 2564 5764 2592
rect 6638 2564 6644 2576
rect 3605 2527 3663 2533
rect 3988 2536 5212 2564
rect 5612 2536 5764 2564
rect 5828 2536 6644 2564
rect 1857 2499 1915 2505
rect 1857 2465 1869 2499
rect 1903 2496 1915 2499
rect 2222 2496 2228 2508
rect 1903 2468 2228 2496
rect 1903 2465 1915 2468
rect 1857 2459 1915 2465
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 2866 2456 2872 2508
rect 2924 2496 2930 2508
rect 2924 2468 3280 2496
rect 2924 2456 2930 2468
rect 3252 2440 3280 2468
rect 3234 2388 3240 2440
rect 3292 2388 3298 2440
rect 3418 2388 3424 2440
rect 3476 2388 3482 2440
rect 2133 2363 2191 2369
rect 2133 2329 2145 2363
rect 2179 2329 2191 2363
rect 2133 2323 2191 2329
rect 2148 2292 2176 2323
rect 2314 2292 2320 2304
rect 2148 2264 2320 2292
rect 2314 2252 2320 2264
rect 2372 2252 2378 2304
rect 3436 2292 3464 2388
rect 3620 2360 3648 2527
rect 3988 2437 4016 2536
rect 4157 2499 4215 2505
rect 4157 2465 4169 2499
rect 4203 2496 4215 2499
rect 4246 2496 4252 2508
rect 4203 2468 4252 2496
rect 4203 2465 4215 2468
rect 4157 2459 4215 2465
rect 4246 2456 4252 2468
rect 4304 2456 4310 2508
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 4341 2431 4399 2437
rect 4341 2428 4353 2431
rect 4120 2400 4353 2428
rect 4120 2388 4126 2400
rect 4341 2397 4353 2400
rect 4387 2397 4399 2431
rect 4341 2391 4399 2397
rect 4798 2388 4804 2440
rect 4856 2388 4862 2440
rect 5612 2437 5640 2536
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 5828 2496 5856 2536
rect 6638 2524 6644 2536
rect 6696 2564 6702 2576
rect 7668 2564 7696 2592
rect 6696 2536 7696 2564
rect 6696 2524 6702 2536
rect 5767 2468 5856 2496
rect 5920 2468 6500 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 5597 2431 5655 2437
rect 5597 2397 5609 2431
rect 5643 2397 5655 2431
rect 5597 2391 5655 2397
rect 4614 2360 4620 2372
rect 3620 2332 4620 2360
rect 4614 2320 4620 2332
rect 4672 2320 4678 2372
rect 4709 2363 4767 2369
rect 4709 2329 4721 2363
rect 4755 2360 4767 2363
rect 4982 2360 4988 2372
rect 4755 2332 4988 2360
rect 4755 2329 4767 2332
rect 4709 2323 4767 2329
rect 4982 2320 4988 2332
rect 5040 2320 5046 2372
rect 5184 2360 5212 2391
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 5920 2428 5948 2468
rect 5868 2400 5948 2428
rect 6472 2428 6500 2468
rect 6822 2428 6828 2440
rect 6472 2400 6828 2428
rect 5868 2388 5874 2400
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 6972 2400 7021 2428
rect 6972 2388 6978 2400
rect 7009 2397 7021 2400
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 6362 2360 6368 2372
rect 5184 2332 6368 2360
rect 6362 2320 6368 2332
rect 6420 2320 6426 2372
rect 6457 2363 6515 2369
rect 6457 2329 6469 2363
rect 6503 2329 6515 2363
rect 6457 2323 6515 2329
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 3436 2264 5365 2292
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 5353 2255 5411 2261
rect 5442 2252 5448 2304
rect 5500 2292 5506 2304
rect 6472 2292 6500 2323
rect 5500 2264 6500 2292
rect 5500 2252 5506 2264
rect 6822 2252 6828 2304
rect 6880 2292 6886 2304
rect 7101 2295 7159 2301
rect 7101 2292 7113 2295
rect 6880 2264 7113 2292
rect 6880 2252 6886 2264
rect 7101 2261 7113 2264
rect 7147 2261 7159 2295
rect 7101 2255 7159 2261
rect 1104 2202 8096 2224
rect 1104 2150 2483 2202
rect 2535 2150 2547 2202
rect 2599 2150 2611 2202
rect 2663 2150 2675 2202
rect 2727 2150 2739 2202
rect 2791 2150 4230 2202
rect 4282 2150 4294 2202
rect 4346 2150 4358 2202
rect 4410 2150 4422 2202
rect 4474 2150 4486 2202
rect 4538 2150 5977 2202
rect 6029 2150 6041 2202
rect 6093 2150 6105 2202
rect 6157 2150 6169 2202
rect 6221 2150 6233 2202
rect 6285 2150 7724 2202
rect 7776 2150 7788 2202
rect 7840 2150 7852 2202
rect 7904 2150 7916 2202
rect 7968 2150 7980 2202
rect 8032 2150 8096 2202
rect 1104 2128 8096 2150
rect 3234 1980 3240 2032
rect 3292 2020 3298 2032
rect 4798 2020 4804 2032
rect 3292 1992 4804 2020
rect 3292 1980 3298 1992
rect 4798 1980 4804 1992
rect 4856 1980 4862 2032
<< via1 >>
rect 2780 8848 2832 8900
rect 2964 8848 3016 8900
rect 4620 8780 4672 8832
rect 5264 8780 5316 8832
rect 2483 8678 2535 8730
rect 2547 8678 2599 8730
rect 2611 8678 2663 8730
rect 2675 8678 2727 8730
rect 2739 8678 2791 8730
rect 4230 8678 4282 8730
rect 4294 8678 4346 8730
rect 4358 8678 4410 8730
rect 4422 8678 4474 8730
rect 4486 8678 4538 8730
rect 5977 8678 6029 8730
rect 6041 8678 6093 8730
rect 6105 8678 6157 8730
rect 6169 8678 6221 8730
rect 6233 8678 6285 8730
rect 7724 8678 7776 8730
rect 7788 8678 7840 8730
rect 7852 8678 7904 8730
rect 7916 8678 7968 8730
rect 7980 8678 8032 8730
rect 2964 8619 3016 8628
rect 2964 8585 2973 8619
rect 2973 8585 3007 8619
rect 3007 8585 3016 8619
rect 2964 8576 3016 8585
rect 2872 8508 2924 8560
rect 1676 8440 1728 8492
rect 2228 8440 2280 8492
rect 3056 8483 3108 8492
rect 3056 8449 3065 8483
rect 3065 8449 3099 8483
rect 3099 8449 3108 8483
rect 3056 8440 3108 8449
rect 3976 8576 4028 8628
rect 5540 8576 5592 8628
rect 5816 8576 5868 8628
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 9036 8576 9088 8628
rect 5264 8508 5316 8560
rect 6368 8508 6420 8560
rect 4160 8440 4212 8492
rect 3884 8372 3936 8424
rect 4620 8440 4672 8492
rect 4988 8440 5040 8492
rect 5080 8440 5132 8492
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 5724 8440 5776 8492
rect 6828 8440 6880 8492
rect 7564 8440 7616 8492
rect 6552 8372 6604 8424
rect 664 8236 716 8288
rect 3148 8304 3200 8356
rect 6276 8304 6328 8356
rect 2504 8236 2556 8288
rect 5172 8279 5224 8288
rect 5172 8245 5181 8279
rect 5181 8245 5215 8279
rect 5215 8245 5224 8279
rect 5172 8236 5224 8245
rect 1823 8134 1875 8186
rect 1887 8134 1939 8186
rect 1951 8134 2003 8186
rect 2015 8134 2067 8186
rect 2079 8134 2131 8186
rect 3570 8134 3622 8186
rect 3634 8134 3686 8186
rect 3698 8134 3750 8186
rect 3762 8134 3814 8186
rect 3826 8134 3878 8186
rect 5317 8134 5369 8186
rect 5381 8134 5433 8186
rect 5445 8134 5497 8186
rect 5509 8134 5561 8186
rect 5573 8134 5625 8186
rect 7064 8134 7116 8186
rect 7128 8134 7180 8186
rect 7192 8134 7244 8186
rect 7256 8134 7308 8186
rect 7320 8134 7372 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 2228 8032 2280 8084
rect 2412 8032 2464 8084
rect 1676 7828 1728 7880
rect 2504 7896 2556 7948
rect 4804 7964 4856 8016
rect 6276 8032 6328 8084
rect 6828 8075 6880 8084
rect 6828 8041 6837 8075
rect 6837 8041 6871 8075
rect 6871 8041 6880 8075
rect 6828 8032 6880 8041
rect 2228 7828 2280 7880
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 2688 7828 2740 7880
rect 6920 7896 6972 7948
rect 1492 7760 1544 7812
rect 1768 7803 1820 7812
rect 1768 7769 1777 7803
rect 1777 7769 1811 7803
rect 1811 7769 1820 7803
rect 1768 7760 1820 7769
rect 2872 7760 2924 7812
rect 2320 7692 2372 7744
rect 4160 7828 4212 7880
rect 4620 7828 4672 7880
rect 4712 7828 4764 7880
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 3332 7692 3384 7744
rect 6460 7803 6512 7812
rect 6460 7769 6469 7803
rect 6469 7769 6503 7803
rect 6503 7769 6512 7803
rect 6460 7760 6512 7769
rect 7104 7803 7156 7812
rect 7104 7769 7113 7803
rect 7113 7769 7147 7803
rect 7147 7769 7156 7803
rect 7104 7760 7156 7769
rect 8208 7828 8260 7880
rect 5540 7692 5592 7744
rect 5816 7692 5868 7744
rect 8116 7692 8168 7744
rect 2483 7590 2535 7642
rect 2547 7590 2599 7642
rect 2611 7590 2663 7642
rect 2675 7590 2727 7642
rect 2739 7590 2791 7642
rect 4230 7590 4282 7642
rect 4294 7590 4346 7642
rect 4358 7590 4410 7642
rect 4422 7590 4474 7642
rect 4486 7590 4538 7642
rect 5977 7590 6029 7642
rect 6041 7590 6093 7642
rect 6105 7590 6157 7642
rect 6169 7590 6221 7642
rect 6233 7590 6285 7642
rect 7724 7590 7776 7642
rect 7788 7590 7840 7642
rect 7852 7590 7904 7642
rect 7916 7590 7968 7642
rect 7980 7590 8032 7642
rect 1768 7488 1820 7540
rect 2412 7488 2464 7540
rect 4160 7488 4212 7540
rect 5172 7488 5224 7540
rect 6460 7488 6512 7540
rect 6552 7488 6604 7540
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 1676 7352 1728 7404
rect 2320 7352 2372 7404
rect 3700 7420 3752 7472
rect 4712 7420 4764 7472
rect 2504 7284 2556 7336
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 5540 7420 5592 7472
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 5816 7352 5868 7404
rect 6368 7352 6420 7404
rect 6552 7352 6604 7404
rect 6644 7352 6696 7404
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 7012 7352 7064 7404
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 3240 7284 3292 7336
rect 3700 7284 3752 7336
rect 4988 7284 5040 7336
rect 5172 7284 5224 7336
rect 7472 7395 7524 7404
rect 7472 7361 7481 7395
rect 7481 7361 7515 7395
rect 7515 7361 7524 7395
rect 7472 7352 7524 7361
rect 5724 7216 5776 7268
rect 3976 7148 4028 7200
rect 5908 7148 5960 7200
rect 6460 7148 6512 7200
rect 7104 7148 7156 7200
rect 1823 7046 1875 7098
rect 1887 7046 1939 7098
rect 1951 7046 2003 7098
rect 2015 7046 2067 7098
rect 2079 7046 2131 7098
rect 3570 7046 3622 7098
rect 3634 7046 3686 7098
rect 3698 7046 3750 7098
rect 3762 7046 3814 7098
rect 3826 7046 3878 7098
rect 5317 7046 5369 7098
rect 5381 7046 5433 7098
rect 5445 7046 5497 7098
rect 5509 7046 5561 7098
rect 5573 7046 5625 7098
rect 7064 7046 7116 7098
rect 7128 7046 7180 7098
rect 7192 7046 7244 7098
rect 7256 7046 7308 7098
rect 7320 7046 7372 7098
rect 940 6808 992 6860
rect 1584 6876 1636 6928
rect 1768 6944 1820 6996
rect 2320 6944 2372 6996
rect 5816 6944 5868 6996
rect 2412 6740 2464 6792
rect 2504 6783 2556 6792
rect 2504 6749 2533 6783
rect 2533 6749 2556 6783
rect 3148 6876 3200 6928
rect 2688 6808 2740 6860
rect 3424 6808 3476 6860
rect 3516 6808 3568 6860
rect 2504 6740 2556 6749
rect 2964 6740 3016 6792
rect 5356 6808 5408 6860
rect 1492 6604 1544 6656
rect 4896 6740 4948 6792
rect 5080 6672 5132 6724
rect 6644 6808 6696 6860
rect 6736 6808 6788 6860
rect 7472 6808 7524 6860
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 3976 6604 4028 6656
rect 4988 6604 5040 6656
rect 5632 6604 5684 6656
rect 5816 6604 5868 6656
rect 7196 6672 7248 6724
rect 2483 6502 2535 6554
rect 2547 6502 2599 6554
rect 2611 6502 2663 6554
rect 2675 6502 2727 6554
rect 2739 6502 2791 6554
rect 4230 6502 4282 6554
rect 4294 6502 4346 6554
rect 4358 6502 4410 6554
rect 4422 6502 4474 6554
rect 4486 6502 4538 6554
rect 5977 6502 6029 6554
rect 6041 6502 6093 6554
rect 6105 6502 6157 6554
rect 6169 6502 6221 6554
rect 6233 6502 6285 6554
rect 7724 6502 7776 6554
rect 7788 6502 7840 6554
rect 7852 6502 7904 6554
rect 7916 6502 7968 6554
rect 7980 6502 8032 6554
rect 1400 6443 1452 6452
rect 1400 6409 1409 6443
rect 1409 6409 1443 6443
rect 1443 6409 1452 6443
rect 1400 6400 1452 6409
rect 2872 6400 2924 6452
rect 3516 6400 3568 6452
rect 3976 6400 4028 6452
rect 3240 6332 3292 6384
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 2228 6239 2280 6248
rect 2228 6205 2237 6239
rect 2237 6205 2271 6239
rect 2271 6205 2280 6239
rect 2228 6196 2280 6205
rect 2780 6196 2832 6248
rect 4068 6332 4120 6384
rect 4712 6332 4764 6384
rect 7104 6332 7156 6384
rect 7380 6375 7432 6384
rect 7380 6341 7389 6375
rect 7389 6341 7423 6375
rect 7423 6341 7432 6375
rect 7380 6332 7432 6341
rect 5356 6264 5408 6316
rect 4068 6239 4120 6248
rect 4068 6205 4077 6239
rect 4077 6205 4111 6239
rect 4111 6205 4120 6239
rect 4068 6196 4120 6205
rect 4620 6196 4672 6248
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 6460 6264 6512 6316
rect 1308 6128 1360 6180
rect 3056 6128 3108 6180
rect 2228 6060 2280 6112
rect 3332 6060 3384 6112
rect 6644 6128 6696 6180
rect 6828 6264 6880 6316
rect 7104 6196 7156 6248
rect 8208 6196 8260 6248
rect 6828 6128 6880 6180
rect 7840 6128 7892 6180
rect 5172 6060 5224 6112
rect 6184 6060 6236 6112
rect 7012 6103 7064 6112
rect 7012 6069 7021 6103
rect 7021 6069 7055 6103
rect 7055 6069 7064 6103
rect 7012 6060 7064 6069
rect 7196 6060 7248 6112
rect 7748 6060 7800 6112
rect 1823 5958 1875 6010
rect 1887 5958 1939 6010
rect 1951 5958 2003 6010
rect 2015 5958 2067 6010
rect 2079 5958 2131 6010
rect 3570 5958 3622 6010
rect 3634 5958 3686 6010
rect 3698 5958 3750 6010
rect 3762 5958 3814 6010
rect 3826 5958 3878 6010
rect 5317 5958 5369 6010
rect 5381 5958 5433 6010
rect 5445 5958 5497 6010
rect 5509 5958 5561 6010
rect 5573 5958 5625 6010
rect 7064 5958 7116 6010
rect 7128 5958 7180 6010
rect 7192 5958 7244 6010
rect 7256 5958 7308 6010
rect 7320 5958 7372 6010
rect 1216 5856 1268 5908
rect 1308 5788 1360 5840
rect 1584 5720 1636 5772
rect 1676 5652 1728 5704
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 2872 5788 2924 5840
rect 2596 5720 2648 5772
rect 1308 5584 1360 5636
rect 3056 5695 3108 5704
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 4068 5856 4120 5908
rect 4988 5856 5040 5908
rect 6460 5856 6512 5908
rect 8116 5856 8168 5908
rect 7380 5788 7432 5840
rect 7748 5788 7800 5840
rect 6644 5720 6696 5772
rect 3976 5652 4028 5704
rect 7840 5652 7892 5704
rect 1676 5516 1728 5568
rect 2044 5516 2096 5568
rect 2412 5516 2464 5568
rect 4160 5584 4212 5636
rect 4712 5584 4764 5636
rect 5908 5627 5960 5636
rect 5908 5593 5917 5627
rect 5917 5593 5951 5627
rect 5951 5593 5960 5627
rect 5908 5584 5960 5593
rect 3240 5516 3292 5568
rect 5172 5516 5224 5568
rect 6184 5516 6236 5568
rect 6644 5516 6696 5568
rect 6828 5516 6880 5568
rect 2483 5414 2535 5466
rect 2547 5414 2599 5466
rect 2611 5414 2663 5466
rect 2675 5414 2727 5466
rect 2739 5414 2791 5466
rect 4230 5414 4282 5466
rect 4294 5414 4346 5466
rect 4358 5414 4410 5466
rect 4422 5414 4474 5466
rect 4486 5414 4538 5466
rect 5977 5414 6029 5466
rect 6041 5414 6093 5466
rect 6105 5414 6157 5466
rect 6169 5414 6221 5466
rect 6233 5414 6285 5466
rect 7724 5414 7776 5466
rect 7788 5414 7840 5466
rect 7852 5414 7904 5466
rect 7916 5414 7968 5466
rect 7980 5414 8032 5466
rect 2228 5312 2280 5364
rect 2044 5244 2096 5296
rect 3976 5312 4028 5364
rect 6368 5312 6420 5364
rect 7472 5312 7524 5364
rect 1584 5176 1636 5228
rect 1308 5108 1360 5160
rect 2504 5219 2556 5228
rect 2504 5185 2513 5219
rect 2513 5185 2547 5219
rect 2547 5185 2556 5219
rect 2504 5176 2556 5185
rect 2780 5219 2832 5228
rect 2780 5185 2789 5219
rect 2789 5185 2823 5219
rect 2823 5185 2832 5219
rect 2780 5176 2832 5185
rect 3332 5176 3384 5228
rect 7656 5244 7708 5296
rect 3056 5108 3108 5160
rect 2504 5040 2556 5092
rect 3148 5083 3200 5092
rect 3148 5049 3157 5083
rect 3157 5049 3191 5083
rect 3191 5049 3200 5083
rect 3148 5040 3200 5049
rect 940 4972 992 5024
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 3056 4972 3108 5024
rect 5908 5040 5960 5092
rect 7380 5219 7432 5228
rect 7380 5185 7389 5219
rect 7389 5185 7423 5219
rect 7423 5185 7432 5219
rect 7380 5176 7432 5185
rect 8116 5176 8168 5228
rect 4160 4972 4212 5024
rect 4620 4972 4672 5024
rect 5816 4972 5868 5024
rect 7656 4972 7708 5024
rect 1823 4870 1875 4922
rect 1887 4870 1939 4922
rect 1951 4870 2003 4922
rect 2015 4870 2067 4922
rect 2079 4870 2131 4922
rect 3570 4870 3622 4922
rect 3634 4870 3686 4922
rect 3698 4870 3750 4922
rect 3762 4870 3814 4922
rect 3826 4870 3878 4922
rect 5317 4870 5369 4922
rect 5381 4870 5433 4922
rect 5445 4870 5497 4922
rect 5509 4870 5561 4922
rect 5573 4870 5625 4922
rect 7064 4870 7116 4922
rect 7128 4870 7180 4922
rect 7192 4870 7244 4922
rect 7256 4870 7308 4922
rect 7320 4870 7372 4922
rect 3056 4768 3108 4820
rect 4896 4768 4948 4820
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 2872 4700 2924 4752
rect 2228 4632 2280 4684
rect 1676 4564 1728 4616
rect 1400 4539 1452 4548
rect 1400 4505 1409 4539
rect 1409 4505 1443 4539
rect 1443 4505 1452 4539
rect 1400 4496 1452 4505
rect 1952 4539 2004 4548
rect 1952 4505 1961 4539
rect 1961 4505 1995 4539
rect 1995 4505 2004 4539
rect 1952 4496 2004 4505
rect 2044 4496 2096 4548
rect 3240 4564 3292 4616
rect 4160 4700 4212 4752
rect 3976 4675 4028 4684
rect 3976 4641 3985 4675
rect 3985 4641 4019 4675
rect 4019 4641 4028 4675
rect 3976 4632 4028 4641
rect 6368 4632 6420 4684
rect 6828 4632 6880 4684
rect 7472 4632 7524 4684
rect 4528 4564 4580 4616
rect 4620 4496 4672 4548
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 3884 4428 3936 4480
rect 4160 4428 4212 4480
rect 8392 4496 8444 4548
rect 5816 4428 5868 4480
rect 2483 4326 2535 4378
rect 2547 4326 2599 4378
rect 2611 4326 2663 4378
rect 2675 4326 2727 4378
rect 2739 4326 2791 4378
rect 4230 4326 4282 4378
rect 4294 4326 4346 4378
rect 4358 4326 4410 4378
rect 4422 4326 4474 4378
rect 4486 4326 4538 4378
rect 5977 4326 6029 4378
rect 6041 4326 6093 4378
rect 6105 4326 6157 4378
rect 6169 4326 6221 4378
rect 6233 4326 6285 4378
rect 7724 4326 7776 4378
rect 7788 4326 7840 4378
rect 7852 4326 7904 4378
rect 7916 4326 7968 4378
rect 7980 4326 8032 4378
rect 1308 4224 1360 4276
rect 1584 4224 1636 4276
rect 3424 4224 3476 4276
rect 1216 4088 1268 4140
rect 1584 4020 1636 4072
rect 1676 4020 1728 4072
rect 2044 4088 2096 4140
rect 4252 4156 4304 4208
rect 5632 4224 5684 4276
rect 5908 4224 5960 4276
rect 5172 4156 5224 4208
rect 2228 4020 2280 4072
rect 2780 4063 2832 4072
rect 2780 4029 2789 4063
rect 2789 4029 2823 4063
rect 2823 4029 2832 4063
rect 2780 4020 2832 4029
rect 6368 4267 6420 4276
rect 6368 4233 6377 4267
rect 6377 4233 6411 4267
rect 6411 4233 6420 4267
rect 6368 4224 6420 4233
rect 7472 4224 7524 4276
rect 7564 4224 7616 4276
rect 7380 4199 7432 4208
rect 7380 4165 7389 4199
rect 7389 4165 7423 4199
rect 7423 4165 7432 4199
rect 7380 4156 7432 4165
rect 8208 4156 8260 4208
rect 2964 4020 3016 4072
rect 6460 4020 6512 4072
rect 6828 4020 6880 4072
rect 7748 4088 7800 4140
rect 7840 4020 7892 4072
rect 20 3884 72 3936
rect 1952 3884 2004 3936
rect 3332 3884 3384 3936
rect 3884 3884 3936 3936
rect 5080 3884 5132 3936
rect 6460 3884 6512 3936
rect 7656 3884 7708 3936
rect 1823 3782 1875 3834
rect 1887 3782 1939 3834
rect 1951 3782 2003 3834
rect 2015 3782 2067 3834
rect 2079 3782 2131 3834
rect 3570 3782 3622 3834
rect 3634 3782 3686 3834
rect 3698 3782 3750 3834
rect 3762 3782 3814 3834
rect 3826 3782 3878 3834
rect 5317 3782 5369 3834
rect 5381 3782 5433 3834
rect 5445 3782 5497 3834
rect 5509 3782 5561 3834
rect 5573 3782 5625 3834
rect 7064 3782 7116 3834
rect 7128 3782 7180 3834
rect 7192 3782 7244 3834
rect 7256 3782 7308 3834
rect 7320 3782 7372 3834
rect 1492 3680 1544 3732
rect 6368 3680 6420 3732
rect 7564 3680 7616 3732
rect 2228 3544 2280 3596
rect 2872 3544 2924 3596
rect 4252 3544 4304 3596
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 4068 3476 4120 3528
rect 5172 3544 5224 3596
rect 6736 3544 6788 3596
rect 2412 3408 2464 3460
rect 5816 3408 5868 3460
rect 5908 3408 5960 3460
rect 6460 3408 6512 3460
rect 7472 3408 7524 3460
rect 7748 3408 7800 3460
rect 7840 3408 7892 3460
rect 3148 3340 3200 3392
rect 3608 3383 3660 3392
rect 3608 3349 3617 3383
rect 3617 3349 3651 3383
rect 3651 3349 3660 3383
rect 3608 3340 3660 3349
rect 3976 3383 4028 3392
rect 3976 3349 3985 3383
rect 3985 3349 4019 3383
rect 4019 3349 4028 3383
rect 3976 3340 4028 3349
rect 5264 3340 5316 3392
rect 7104 3340 7156 3392
rect 2483 3238 2535 3290
rect 2547 3238 2599 3290
rect 2611 3238 2663 3290
rect 2675 3238 2727 3290
rect 2739 3238 2791 3290
rect 4230 3238 4282 3290
rect 4294 3238 4346 3290
rect 4358 3238 4410 3290
rect 4422 3238 4474 3290
rect 4486 3238 4538 3290
rect 5977 3238 6029 3290
rect 6041 3238 6093 3290
rect 6105 3238 6157 3290
rect 6169 3238 6221 3290
rect 6233 3238 6285 3290
rect 7724 3238 7776 3290
rect 7788 3238 7840 3290
rect 7852 3238 7904 3290
rect 7916 3238 7968 3290
rect 7980 3238 8032 3290
rect 1676 3136 1728 3188
rect 2412 3136 2464 3188
rect 3424 3136 3476 3188
rect 4712 3136 4764 3188
rect 5908 3179 5960 3188
rect 5908 3145 5917 3179
rect 5917 3145 5951 3179
rect 5951 3145 5960 3179
rect 5908 3136 5960 3145
rect 6368 3136 6420 3188
rect 7472 3136 7524 3188
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 1584 2932 1636 2984
rect 2228 2932 2280 2984
rect 4160 3068 4212 3120
rect 4620 3068 4672 3120
rect 6552 3111 6604 3120
rect 6552 3077 6561 3111
rect 6561 3077 6595 3111
rect 6595 3077 6604 3111
rect 6552 3068 6604 3077
rect 6828 3068 6880 3120
rect 5264 3043 5316 3052
rect 5264 3009 5273 3043
rect 5273 3009 5307 3043
rect 5307 3009 5316 3043
rect 5264 3000 5316 3009
rect 5724 3000 5776 3052
rect 3424 2932 3476 2984
rect 3608 2932 3660 2984
rect 4988 2975 5040 2984
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 5172 2932 5224 2984
rect 7104 3000 7156 3052
rect 7564 3068 7616 3120
rect 2688 2864 2740 2916
rect 4252 2864 4304 2916
rect 4160 2796 4212 2848
rect 6828 2796 6880 2848
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 1823 2694 1875 2746
rect 1887 2694 1939 2746
rect 1951 2694 2003 2746
rect 2015 2694 2067 2746
rect 2079 2694 2131 2746
rect 3570 2694 3622 2746
rect 3634 2694 3686 2746
rect 3698 2694 3750 2746
rect 3762 2694 3814 2746
rect 3826 2694 3878 2746
rect 5317 2694 5369 2746
rect 5381 2694 5433 2746
rect 5445 2694 5497 2746
rect 5509 2694 5561 2746
rect 5573 2694 5625 2746
rect 7064 2694 7116 2746
rect 7128 2694 7180 2746
rect 7192 2694 7244 2746
rect 7256 2694 7308 2746
rect 7320 2694 7372 2746
rect 3976 2592 4028 2644
rect 5172 2592 5224 2644
rect 5724 2592 5776 2644
rect 7656 2592 7708 2644
rect 2228 2456 2280 2508
rect 2872 2456 2924 2508
rect 3240 2388 3292 2440
rect 3424 2388 3476 2440
rect 2320 2252 2372 2304
rect 4252 2456 4304 2508
rect 4068 2388 4120 2440
rect 4804 2431 4856 2440
rect 4804 2397 4813 2431
rect 4813 2397 4847 2431
rect 4847 2397 4856 2431
rect 4804 2388 4856 2397
rect 6644 2524 6696 2576
rect 4620 2320 4672 2372
rect 4988 2320 5040 2372
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 6828 2431 6880 2440
rect 5816 2388 5868 2397
rect 6828 2397 6837 2431
rect 6837 2397 6871 2431
rect 6871 2397 6880 2431
rect 6828 2388 6880 2397
rect 6920 2388 6972 2440
rect 6368 2320 6420 2372
rect 5448 2252 5500 2304
rect 6828 2252 6880 2304
rect 2483 2150 2535 2202
rect 2547 2150 2599 2202
rect 2611 2150 2663 2202
rect 2675 2150 2727 2202
rect 2739 2150 2791 2202
rect 4230 2150 4282 2202
rect 4294 2150 4346 2202
rect 4358 2150 4410 2202
rect 4422 2150 4474 2202
rect 4486 2150 4538 2202
rect 5977 2150 6029 2202
rect 6041 2150 6093 2202
rect 6105 2150 6157 2202
rect 6169 2150 6221 2202
rect 6233 2150 6285 2202
rect 7724 2150 7776 2202
rect 7788 2150 7840 2202
rect 7852 2150 7904 2202
rect 7916 2150 7968 2202
rect 7980 2150 8032 2202
rect 3240 1980 3292 2032
rect 4804 1980 4856 2032
<< metal2 >>
rect 662 10548 718 11348
rect 2594 10690 2650 11348
rect 2594 10662 2728 10690
rect 2594 10548 2650 10662
rect 676 8294 704 10548
rect 2700 9466 2728 10662
rect 3882 10548 3938 11348
rect 5814 10548 5870 11348
rect 7746 10548 7802 11348
rect 9034 10548 9090 11348
rect 2778 10296 2834 10305
rect 2834 10254 2912 10282
rect 2778 10231 2834 10240
rect 2700 9438 2820 9466
rect 1490 8936 1546 8945
rect 2792 8906 2820 9438
rect 1490 8871 1546 8880
rect 2780 8900 2832 8906
rect 664 8288 716 8294
rect 664 8230 716 8236
rect 1504 8090 1532 8871
rect 2780 8842 2832 8848
rect 2483 8732 2791 8741
rect 2483 8730 2489 8732
rect 2545 8730 2569 8732
rect 2625 8730 2649 8732
rect 2705 8730 2729 8732
rect 2785 8730 2791 8732
rect 2545 8678 2547 8730
rect 2727 8678 2729 8730
rect 2483 8676 2489 8678
rect 2545 8676 2569 8678
rect 2625 8676 2649 8678
rect 2705 8676 2729 8678
rect 2785 8676 2791 8678
rect 2483 8667 2791 8676
rect 2884 8566 2912 10254
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 2976 8634 3004 8842
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1688 7886 1716 8434
rect 1823 8188 2131 8197
rect 1823 8186 1829 8188
rect 1885 8186 1909 8188
rect 1965 8186 1989 8188
rect 2045 8186 2069 8188
rect 2125 8186 2131 8188
rect 1885 8134 1887 8186
rect 2067 8134 2069 8186
rect 1823 8132 1829 8134
rect 1885 8132 1909 8134
rect 1965 8132 1989 8134
rect 2045 8132 2069 8134
rect 2125 8132 2131 8134
rect 1823 8123 2131 8132
rect 2240 8090 2268 8434
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2424 7886 2452 8026
rect 2516 7954 2544 8230
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2412 7880 2464 7886
rect 2688 7880 2740 7886
rect 2412 7822 2464 7828
rect 2686 7848 2688 7857
rect 2740 7848 2742 7857
rect 1492 7812 1544 7818
rect 1492 7754 1544 7760
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 938 6896 994 6905
rect 938 6831 940 6840
rect 992 6831 994 6840
rect 940 6802 992 6808
rect 1214 6760 1270 6769
rect 1214 6695 1270 6704
rect 1228 5914 1256 6695
rect 1412 6458 1440 7346
rect 1504 6780 1532 7754
rect 1780 7546 1808 7754
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6934 1624 7142
rect 1584 6928 1636 6934
rect 1584 6870 1636 6876
rect 1504 6752 1624 6780
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1308 6180 1360 6186
rect 1308 6122 1360 6128
rect 1216 5908 1268 5914
rect 1216 5850 1268 5856
rect 940 5024 992 5030
rect 940 4966 992 4972
rect 952 4865 980 4966
rect 938 4856 994 4865
rect 938 4791 994 4800
rect 1228 4146 1256 5850
rect 1320 5846 1348 6122
rect 1308 5840 1360 5846
rect 1308 5782 1360 5788
rect 1308 5636 1360 5642
rect 1308 5578 1360 5584
rect 1320 5166 1348 5578
rect 1308 5160 1360 5166
rect 1308 5102 1360 5108
rect 1320 4282 1348 5102
rect 1400 4548 1452 4554
rect 1400 4490 1452 4496
rect 1308 4276 1360 4282
rect 1308 4218 1360 4224
rect 1216 4140 1268 4146
rect 1216 4082 1268 4088
rect 20 3936 72 3942
rect 20 3878 72 3884
rect 32 800 60 3878
rect 1412 2774 1440 4490
rect 1504 3738 1532 6598
rect 1596 5778 1624 6752
rect 1688 6322 1716 7346
rect 1823 7100 2131 7109
rect 1823 7098 1829 7100
rect 1885 7098 1909 7100
rect 1965 7098 1989 7100
rect 2045 7098 2069 7100
rect 2125 7098 2131 7100
rect 1885 7046 1887 7098
rect 2067 7046 2069 7098
rect 1823 7044 1829 7046
rect 1885 7044 1909 7046
rect 1965 7044 1989 7046
rect 2045 7044 2069 7046
rect 2125 7044 2131 7046
rect 1823 7035 2131 7044
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1780 6100 1808 6938
rect 2240 6882 2268 7822
rect 2686 7783 2742 7792
rect 2872 7812 2924 7818
rect 2872 7754 2924 7760
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2332 7410 2360 7686
rect 2483 7644 2791 7653
rect 2483 7642 2489 7644
rect 2545 7642 2569 7644
rect 2625 7642 2649 7644
rect 2705 7642 2729 7644
rect 2785 7642 2791 7644
rect 2545 7590 2547 7642
rect 2727 7590 2729 7642
rect 2483 7588 2489 7590
rect 2545 7588 2569 7590
rect 2625 7588 2649 7590
rect 2705 7588 2729 7590
rect 2785 7588 2791 7590
rect 2483 7579 2791 7588
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2332 7002 2360 7346
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2240 6854 2360 6882
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2240 6361 2268 6598
rect 2226 6352 2282 6361
rect 2226 6287 2282 6296
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2240 6118 2268 6190
rect 1688 6072 1808 6100
rect 2228 6112 2280 6118
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1688 5710 1716 6072
rect 2228 6054 2280 6060
rect 1823 6012 2131 6021
rect 1823 6010 1829 6012
rect 1885 6010 1909 6012
rect 1965 6010 1989 6012
rect 2045 6010 2069 6012
rect 2125 6010 2131 6012
rect 1885 5958 1887 6010
rect 2067 5958 2069 6010
rect 1823 5956 1829 5958
rect 1885 5956 1909 5958
rect 1965 5956 1989 5958
rect 2045 5956 2069 5958
rect 2125 5956 2131 5958
rect 1823 5947 2131 5956
rect 2332 5896 2360 6854
rect 2424 6798 2452 7482
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2516 6798 2544 7278
rect 2686 7032 2742 7041
rect 2686 6967 2742 6976
rect 2700 6866 2728 6967
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2504 6792 2556 6798
rect 2700 6769 2728 6802
rect 2504 6734 2556 6740
rect 2686 6760 2742 6769
rect 2424 6338 2452 6734
rect 2686 6695 2742 6704
rect 2483 6556 2791 6565
rect 2483 6554 2489 6556
rect 2545 6554 2569 6556
rect 2625 6554 2649 6556
rect 2705 6554 2729 6556
rect 2785 6554 2791 6556
rect 2545 6502 2547 6554
rect 2727 6502 2729 6554
rect 2483 6500 2489 6502
rect 2545 6500 2569 6502
rect 2625 6500 2649 6502
rect 2705 6500 2729 6502
rect 2785 6500 2791 6502
rect 2483 6491 2791 6500
rect 2884 6458 2912 7754
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2976 6474 3004 6734
rect 3068 6662 3096 8434
rect 3896 8430 3924 10548
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4230 8732 4538 8741
rect 4230 8730 4236 8732
rect 4292 8730 4316 8732
rect 4372 8730 4396 8732
rect 4452 8730 4476 8732
rect 4532 8730 4538 8732
rect 4292 8678 4294 8730
rect 4474 8678 4476 8730
rect 4230 8676 4236 8678
rect 4292 8676 4316 8678
rect 4372 8676 4396 8678
rect 4452 8676 4476 8678
rect 4532 8676 4538 8678
rect 4230 8667 4538 8676
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3160 7041 3188 8298
rect 3570 8188 3878 8197
rect 3570 8186 3576 8188
rect 3632 8186 3656 8188
rect 3712 8186 3736 8188
rect 3792 8186 3816 8188
rect 3872 8186 3878 8188
rect 3632 8134 3634 8186
rect 3814 8134 3816 8186
rect 3570 8132 3576 8134
rect 3632 8132 3656 8134
rect 3712 8132 3736 8134
rect 3792 8132 3816 8134
rect 3872 8132 3878 8134
rect 3570 8123 3878 8132
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3146 7032 3202 7041
rect 3146 6967 3202 6976
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2872 6452 2924 6458
rect 2976 6446 3096 6474
rect 2872 6394 2924 6400
rect 2424 6310 2636 6338
rect 2056 5868 2360 5896
rect 2056 5710 2084 5868
rect 2608 5794 2636 6310
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2792 6066 2820 6190
rect 3068 6186 3096 6446
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 2792 6038 3004 6066
rect 2240 5778 2636 5794
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2240 5772 2648 5778
rect 2240 5766 2596 5772
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 4282 1624 5170
rect 1688 4622 1716 5510
rect 2056 5302 2084 5510
rect 2240 5370 2268 5766
rect 2596 5714 2648 5720
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2044 5296 2096 5302
rect 2044 5238 2096 5244
rect 2148 5086 2360 5114
rect 2148 5030 2176 5086
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 1823 4924 2131 4933
rect 1823 4922 1829 4924
rect 1885 4922 1909 4924
rect 1965 4922 1989 4924
rect 2045 4922 2069 4924
rect 2125 4922 2131 4924
rect 1885 4870 1887 4922
rect 2067 4870 2069 4922
rect 1823 4868 1829 4870
rect 1885 4868 1909 4870
rect 1965 4868 1989 4870
rect 2045 4868 2069 4870
rect 2125 4868 2131 4870
rect 1823 4859 2131 4868
rect 2240 4690 2268 4966
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1952 4548 2004 4554
rect 1952 4490 2004 4496
rect 2044 4548 2096 4554
rect 2044 4490 2096 4496
rect 1584 4276 1636 4282
rect 1584 4218 1636 4224
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1492 3732 1544 3738
rect 1492 3674 1544 3680
rect 1596 2990 1624 4014
rect 1688 3194 1716 4014
rect 1964 3942 1992 4490
rect 2056 4146 2084 4490
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1823 3836 2131 3845
rect 1823 3834 1829 3836
rect 1885 3834 1909 3836
rect 1965 3834 1989 3836
rect 2045 3834 2069 3836
rect 2125 3834 2131 3836
rect 1885 3782 1887 3834
rect 2067 3782 2069 3834
rect 1823 3780 1829 3782
rect 1885 3780 1909 3782
rect 1965 3780 1989 3782
rect 2045 3780 2069 3782
rect 2125 3780 2131 3782
rect 1823 3771 2131 3780
rect 2240 3602 2268 4014
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 2056 2938 2084 2994
rect 2240 2990 2268 3538
rect 2228 2984 2280 2990
rect 2134 2952 2190 2961
rect 2056 2910 2134 2938
rect 2228 2926 2280 2932
rect 2134 2887 2190 2896
rect 1320 2746 1440 2774
rect 1823 2748 2131 2757
rect 1823 2746 1829 2748
rect 1885 2746 1909 2748
rect 1965 2746 1989 2748
rect 2045 2746 2069 2748
rect 2125 2746 2131 2748
rect 1320 800 1348 2746
rect 1885 2694 1887 2746
rect 2067 2694 2069 2746
rect 1823 2692 1829 2694
rect 1885 2692 1909 2694
rect 1965 2692 1989 2694
rect 2045 2692 2069 2694
rect 2125 2692 2131 2694
rect 1823 2683 2131 2692
rect 2240 2514 2268 2926
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2332 2310 2360 5086
rect 2424 3466 2452 5510
rect 2483 5468 2791 5477
rect 2483 5466 2489 5468
rect 2545 5466 2569 5468
rect 2625 5466 2649 5468
rect 2705 5466 2729 5468
rect 2785 5466 2791 5468
rect 2545 5414 2547 5466
rect 2727 5414 2729 5466
rect 2483 5412 2489 5414
rect 2545 5412 2569 5414
rect 2625 5412 2649 5414
rect 2705 5412 2729 5414
rect 2785 5412 2791 5414
rect 2483 5403 2791 5412
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2780 5228 2832 5234
rect 2884 5216 2912 5782
rect 2832 5188 2912 5216
rect 2780 5170 2832 5176
rect 2516 5098 2544 5170
rect 2792 5137 2820 5170
rect 2778 5128 2834 5137
rect 2504 5092 2556 5098
rect 2778 5063 2834 5072
rect 2504 5034 2556 5040
rect 2872 4752 2924 4758
rect 2872 4694 2924 4700
rect 2483 4380 2791 4389
rect 2483 4378 2489 4380
rect 2545 4378 2569 4380
rect 2625 4378 2649 4380
rect 2705 4378 2729 4380
rect 2785 4378 2791 4380
rect 2545 4326 2547 4378
rect 2727 4326 2729 4378
rect 2483 4324 2489 4326
rect 2545 4324 2569 4326
rect 2625 4324 2649 4326
rect 2705 4324 2729 4326
rect 2785 4324 2791 4326
rect 2483 4315 2791 4324
rect 2884 4162 2912 4694
rect 2792 4134 2912 4162
rect 2792 4078 2820 4134
rect 2976 4078 3004 6038
rect 3068 5710 3096 6122
rect 3160 5710 3188 6870
rect 3252 6390 3280 7278
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3344 6118 3372 7686
rect 3700 7472 3752 7478
rect 3700 7414 3752 7420
rect 3712 7342 3740 7414
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3988 7206 4016 8570
rect 4632 8498 4660 8774
rect 5276 8566 5304 8774
rect 5828 8634 5856 10548
rect 7102 9616 7158 9625
rect 7102 9551 7158 9560
rect 5977 8732 6285 8741
rect 5977 8730 5983 8732
rect 6039 8730 6063 8732
rect 6119 8730 6143 8732
rect 6199 8730 6223 8732
rect 6279 8730 6285 8732
rect 6039 8678 6041 8730
rect 6221 8678 6223 8730
rect 5977 8676 5983 8678
rect 6039 8676 6063 8678
rect 6119 8676 6143 8678
rect 6199 8676 6223 8678
rect 6279 8676 6285 8678
rect 5977 8667 6285 8676
rect 7116 8634 7144 9551
rect 7760 8922 7788 10548
rect 7668 8894 7788 8922
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4172 7886 4200 8434
rect 4632 7886 4660 8434
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4172 7546 4200 7822
rect 4230 7644 4538 7653
rect 4230 7642 4236 7644
rect 4292 7642 4316 7644
rect 4372 7642 4396 7644
rect 4452 7642 4476 7644
rect 4532 7642 4538 7644
rect 4292 7590 4294 7642
rect 4474 7590 4476 7642
rect 4230 7588 4236 7590
rect 4292 7588 4316 7590
rect 4372 7588 4396 7590
rect 4452 7588 4476 7590
rect 4532 7588 4538 7590
rect 4230 7579 4538 7588
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4724 7478 4752 7822
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3570 7100 3878 7109
rect 3570 7098 3576 7100
rect 3632 7098 3656 7100
rect 3712 7098 3736 7100
rect 3792 7098 3816 7100
rect 3872 7098 3878 7100
rect 3632 7046 3634 7098
rect 3814 7046 3816 7098
rect 3570 7044 3576 7046
rect 3632 7044 3656 7046
rect 3712 7044 3736 7046
rect 3792 7044 3816 7046
rect 3872 7044 3878 7046
rect 3570 7035 3878 7044
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3068 5166 3096 5646
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 3068 4826 3096 4966
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 3160 4298 3188 5034
rect 3252 4622 3280 5510
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3068 4270 3188 4298
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 2483 3292 2791 3301
rect 2483 3290 2489 3292
rect 2545 3290 2569 3292
rect 2625 3290 2649 3292
rect 2705 3290 2729 3292
rect 2785 3290 2791 3292
rect 2545 3238 2547 3290
rect 2727 3238 2729 3290
rect 2483 3236 2489 3238
rect 2545 3236 2569 3238
rect 2625 3236 2649 3238
rect 2705 3236 2729 3238
rect 2785 3236 2791 3238
rect 2483 3227 2791 3236
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2424 3074 2452 3130
rect 2424 3046 2728 3074
rect 2700 2922 2728 3046
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 2884 2514 2912 3538
rect 3068 2774 3096 4270
rect 3252 4026 3280 4422
rect 3160 3998 3280 4026
rect 3160 3398 3188 3998
rect 3344 3942 3372 5170
rect 3436 4468 3464 6802
rect 3528 6458 3556 6802
rect 3988 6662 4016 7142
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3570 6012 3878 6021
rect 3570 6010 3576 6012
rect 3632 6010 3656 6012
rect 3712 6010 3736 6012
rect 3792 6010 3816 6012
rect 3872 6010 3878 6012
rect 3632 5958 3634 6010
rect 3814 5958 3816 6010
rect 3570 5956 3576 5958
rect 3632 5956 3656 5958
rect 3712 5956 3736 5958
rect 3792 5956 3816 5958
rect 3872 5956 3878 5958
rect 3570 5947 3878 5956
rect 3988 5710 4016 6394
rect 4080 6390 4108 7346
rect 4230 6556 4538 6565
rect 4230 6554 4236 6556
rect 4292 6554 4316 6556
rect 4372 6554 4396 6556
rect 4452 6554 4476 6556
rect 4532 6554 4538 6556
rect 4292 6502 4294 6554
rect 4474 6502 4476 6554
rect 4230 6500 4236 6502
rect 4292 6500 4316 6502
rect 4372 6500 4396 6502
rect 4452 6500 4476 6502
rect 4532 6500 4538 6502
rect 4230 6491 4538 6500
rect 4724 6390 4752 7414
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4080 5914 4108 6190
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3988 5370 4016 5646
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4172 5522 4200 5578
rect 4080 5494 4200 5522
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3570 4924 3878 4933
rect 3570 4922 3576 4924
rect 3632 4922 3656 4924
rect 3712 4922 3736 4924
rect 3792 4922 3816 4924
rect 3872 4922 3878 4924
rect 3632 4870 3634 4922
rect 3814 4870 3816 4922
rect 3570 4868 3576 4870
rect 3632 4868 3656 4870
rect 3712 4868 3736 4870
rect 3792 4868 3816 4870
rect 3872 4868 3878 4870
rect 3570 4859 3878 4868
rect 3988 4690 4016 5306
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3884 4480 3936 4486
rect 3436 4440 3556 4468
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3436 3194 3464 4218
rect 3528 4049 3556 4440
rect 3884 4422 3936 4428
rect 3514 4040 3570 4049
rect 3514 3975 3570 3984
rect 3896 3942 3924 4422
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3570 3836 3878 3845
rect 3570 3834 3576 3836
rect 3632 3834 3656 3836
rect 3712 3834 3736 3836
rect 3792 3834 3816 3836
rect 3872 3834 3878 3836
rect 3632 3782 3634 3834
rect 3814 3782 3816 3834
rect 3570 3780 3576 3782
rect 3632 3780 3656 3782
rect 3712 3780 3736 3782
rect 3792 3780 3816 3782
rect 3872 3780 3878 3782
rect 3570 3771 3878 3780
rect 4080 3534 4108 5494
rect 4230 5468 4538 5477
rect 4230 5466 4236 5468
rect 4292 5466 4316 5468
rect 4372 5466 4396 5468
rect 4452 5466 4476 5468
rect 4532 5466 4538 5468
rect 4292 5414 4294 5466
rect 4474 5414 4476 5466
rect 4230 5412 4236 5414
rect 4292 5412 4316 5414
rect 4372 5412 4396 5414
rect 4452 5412 4476 5414
rect 4532 5412 4538 5414
rect 4230 5403 4538 5412
rect 4632 5114 4660 6190
rect 4724 5642 4752 6326
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4540 5086 4752 5114
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4172 4758 4200 4966
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 4540 4622 4568 5086
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4632 4554 4660 4966
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3620 2990 3648 3334
rect 3804 3176 3832 3470
rect 3976 3392 4028 3398
rect 4028 3340 4108 3346
rect 3976 3334 4108 3340
rect 3988 3318 4108 3334
rect 3804 3148 4016 3176
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3068 2746 3188 2774
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2320 2304 2372 2310
rect 2320 2246 2372 2252
rect 2483 2204 2791 2213
rect 2483 2202 2489 2204
rect 2545 2202 2569 2204
rect 2625 2202 2649 2204
rect 2705 2202 2729 2204
rect 2785 2202 2791 2204
rect 2545 2150 2547 2202
rect 2727 2150 2729 2202
rect 2483 2148 2489 2150
rect 2545 2148 2569 2150
rect 2625 2148 2649 2150
rect 2705 2148 2729 2150
rect 2785 2148 2791 2150
rect 2483 2139 2791 2148
rect 3160 1465 3188 2746
rect 3436 2446 3464 2926
rect 3570 2748 3878 2757
rect 3570 2746 3576 2748
rect 3632 2746 3656 2748
rect 3712 2746 3736 2748
rect 3792 2746 3816 2748
rect 3872 2746 3878 2748
rect 3632 2694 3634 2746
rect 3814 2694 3816 2746
rect 3570 2692 3576 2694
rect 3632 2692 3656 2694
rect 3712 2692 3736 2694
rect 3792 2692 3816 2694
rect 3872 2692 3878 2694
rect 3570 2683 3878 2692
rect 3988 2650 4016 3148
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4080 2446 4108 3318
rect 4172 3126 4200 4422
rect 4230 4380 4538 4389
rect 4230 4378 4236 4380
rect 4292 4378 4316 4380
rect 4372 4378 4396 4380
rect 4452 4378 4476 4380
rect 4532 4378 4538 4380
rect 4292 4326 4294 4378
rect 4474 4326 4476 4378
rect 4230 4324 4236 4326
rect 4292 4324 4316 4326
rect 4372 4324 4396 4326
rect 4452 4324 4476 4326
rect 4532 4324 4538 4326
rect 4230 4315 4538 4324
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4264 3602 4292 4150
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4230 3292 4538 3301
rect 4230 3290 4236 3292
rect 4292 3290 4316 3292
rect 4372 3290 4396 3292
rect 4452 3290 4476 3292
rect 4532 3290 4538 3292
rect 4292 3238 4294 3290
rect 4474 3238 4476 3290
rect 4230 3236 4236 3238
rect 4292 3236 4316 3238
rect 4372 3236 4396 3238
rect 4452 3236 4476 3238
rect 4532 3236 4538 3238
rect 4230 3227 4538 3236
rect 4632 3126 4660 4490
rect 4724 3194 4752 5086
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 3252 2038 3280 2382
rect 3240 2032 3292 2038
rect 3240 1974 3292 1980
rect 3146 1456 3202 1465
rect 3146 1391 3202 1400
rect 3252 870 3372 898
rect 3252 800 3280 870
rect 18 0 74 800
rect 1306 0 1362 800
rect 3238 0 3294 800
rect 3344 785 3372 870
rect 4172 785 4200 2790
rect 4264 2514 4292 2858
rect 4724 2774 4752 3130
rect 4632 2746 4752 2774
rect 4816 2774 4844 7958
rect 5000 7342 5028 8434
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 4826 4936 6734
rect 5092 6730 5120 8434
rect 5552 8430 5580 8570
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7546 5212 8230
rect 5317 8188 5625 8197
rect 5317 8186 5323 8188
rect 5379 8186 5403 8188
rect 5459 8186 5483 8188
rect 5539 8186 5563 8188
rect 5619 8186 5625 8188
rect 5379 8134 5381 8186
rect 5561 8134 5563 8186
rect 5317 8132 5323 8134
rect 5379 8132 5403 8134
rect 5459 8132 5483 8134
rect 5539 8132 5563 8134
rect 5619 8132 5625 8134
rect 5317 8123 5625 8132
rect 5262 7848 5318 7857
rect 5262 7783 5318 7792
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5276 7410 5304 7783
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5552 7478 5580 7686
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5000 5914 5028 6598
rect 5184 6118 5212 7278
rect 5736 7274 5764 8434
rect 6276 8356 6328 8362
rect 6276 8298 6328 8304
rect 6288 8090 6316 8298
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5828 7410 5856 7686
rect 5977 7644 6285 7653
rect 5977 7642 5983 7644
rect 6039 7642 6063 7644
rect 6119 7642 6143 7644
rect 6199 7642 6223 7644
rect 6279 7642 6285 7644
rect 6039 7590 6041 7642
rect 6221 7590 6223 7642
rect 5977 7588 5983 7590
rect 6039 7588 6063 7590
rect 6119 7588 6143 7590
rect 6199 7588 6223 7590
rect 6279 7588 6285 7590
rect 5977 7579 6285 7588
rect 6380 7410 6408 8502
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6472 7546 6500 7754
rect 6564 7546 6592 8366
rect 6840 8090 6868 8434
rect 7064 8188 7372 8197
rect 7064 8186 7070 8188
rect 7126 8186 7150 8188
rect 7206 8186 7230 8188
rect 7286 8186 7310 8188
rect 7366 8186 7372 8188
rect 7126 8134 7128 8186
rect 7308 8134 7310 8186
rect 7064 8132 7070 8134
rect 7126 8132 7150 8134
rect 7206 8132 7230 8134
rect 7286 8132 7310 8134
rect 7366 8132 7372 8134
rect 7064 8123 7372 8132
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 5317 7100 5625 7109
rect 5317 7098 5323 7100
rect 5379 7098 5403 7100
rect 5459 7098 5483 7100
rect 5539 7098 5563 7100
rect 5619 7098 5625 7100
rect 5379 7046 5381 7098
rect 5561 7046 5563 7098
rect 5317 7044 5323 7046
rect 5379 7044 5403 7046
rect 5459 7044 5483 7046
rect 5539 7044 5563 7046
rect 5619 7044 5625 7046
rect 5317 7035 5625 7044
rect 5828 7002 5856 7346
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5368 6322 5396 6802
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5172 6112 5224 6118
rect 5644 6100 5672 6598
rect 5644 6072 5764 6100
rect 5172 6054 5224 6060
rect 5317 6012 5625 6021
rect 5317 6010 5323 6012
rect 5379 6010 5403 6012
rect 5459 6010 5483 6012
rect 5539 6010 5563 6012
rect 5619 6010 5625 6012
rect 5379 5958 5381 6010
rect 5561 5958 5563 6010
rect 5317 5956 5323 5958
rect 5379 5956 5403 5958
rect 5459 5956 5483 5958
rect 5539 5956 5563 5958
rect 5619 5956 5625 5958
rect 5317 5947 5625 5956
rect 4988 5908 5040 5914
rect 5040 5868 5120 5896
rect 4988 5850 5040 5856
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5092 4570 5120 5868
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5000 4542 5120 4570
rect 5000 2990 5028 4542
rect 5184 4214 5212 5510
rect 5317 4924 5625 4933
rect 5317 4922 5323 4924
rect 5379 4922 5403 4924
rect 5459 4922 5483 4924
rect 5539 4922 5563 4924
rect 5619 4922 5625 4924
rect 5379 4870 5381 4922
rect 5561 4870 5563 4922
rect 5317 4868 5323 4870
rect 5379 4868 5403 4870
rect 5459 4868 5483 4870
rect 5539 4868 5563 4870
rect 5619 4868 5625 4870
rect 5317 4859 5625 4868
rect 5632 4276 5684 4282
rect 5736 4264 5764 6072
rect 5828 5030 5856 6598
rect 5920 5642 5948 7142
rect 5977 6556 6285 6565
rect 5977 6554 5983 6556
rect 6039 6554 6063 6556
rect 6119 6554 6143 6556
rect 6199 6554 6223 6556
rect 6279 6554 6285 6556
rect 6039 6502 6041 6554
rect 6221 6502 6223 6554
rect 5977 6500 5983 6502
rect 6039 6500 6063 6502
rect 6119 6500 6143 6502
rect 6199 6500 6223 6502
rect 6279 6500 6285 6502
rect 5977 6491 6285 6500
rect 6380 6440 6408 7346
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6196 6412 6408 6440
rect 6196 6118 6224 6412
rect 6472 6322 6500 7142
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6380 6225 6408 6258
rect 6366 6216 6422 6225
rect 6366 6151 6422 6160
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 6196 5574 6224 6054
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 5977 5468 6285 5477
rect 5977 5466 5983 5468
rect 6039 5466 6063 5468
rect 6119 5466 6143 5468
rect 6199 5466 6223 5468
rect 6279 5466 6285 5468
rect 6039 5414 6041 5466
rect 6221 5414 6223 5466
rect 5977 5412 5983 5414
rect 6039 5412 6063 5414
rect 6119 5412 6143 5414
rect 6199 5412 6223 5414
rect 6279 5412 6285 5414
rect 5977 5403 6285 5412
rect 6380 5370 6408 6151
rect 6472 5914 6500 6258
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5684 4236 5764 4264
rect 5632 4218 5684 4224
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 4816 2746 4936 2774
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 4632 2378 4660 2746
rect 4804 2440 4856 2446
rect 4908 2417 4936 2746
rect 4804 2382 4856 2388
rect 4894 2408 4950 2417
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 4230 2204 4538 2213
rect 4230 2202 4236 2204
rect 4292 2202 4316 2204
rect 4372 2202 4396 2204
rect 4452 2202 4476 2204
rect 4532 2202 4538 2204
rect 4292 2150 4294 2202
rect 4474 2150 4476 2202
rect 4230 2148 4236 2150
rect 4292 2148 4316 2150
rect 4372 2148 4396 2150
rect 4452 2148 4476 2150
rect 4532 2148 4538 2150
rect 4230 2139 4538 2148
rect 4816 2038 4844 2382
rect 4894 2343 4950 2352
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 4804 2032 4856 2038
rect 4804 1974 4856 1980
rect 5000 1170 5028 2314
rect 5092 2292 5120 3878
rect 5184 3602 5212 4150
rect 5317 3836 5625 3845
rect 5317 3834 5323 3836
rect 5379 3834 5403 3836
rect 5459 3834 5483 3836
rect 5539 3834 5563 3836
rect 5619 3834 5625 3836
rect 5379 3782 5381 3834
rect 5561 3782 5563 3834
rect 5317 3780 5323 3782
rect 5379 3780 5403 3782
rect 5459 3780 5483 3782
rect 5539 3780 5563 3782
rect 5619 3780 5625 3782
rect 5317 3771 5625 3780
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5828 3466 5856 4422
rect 5920 4282 5948 5034
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 5977 4380 6285 4389
rect 5977 4378 5983 4380
rect 6039 4378 6063 4380
rect 6119 4378 6143 4380
rect 6199 4378 6223 4380
rect 6279 4378 6285 4380
rect 6039 4326 6041 4378
rect 6221 4326 6223 4378
rect 5977 4324 5983 4326
rect 6039 4324 6063 4326
rect 6119 4324 6143 4326
rect 6199 4324 6223 4326
rect 6279 4324 6285 4326
rect 5977 4315 6285 4324
rect 6380 4282 6408 4626
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6472 4078 6500 5850
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5276 3058 5304 3334
rect 5920 3194 5948 3402
rect 5977 3292 6285 3301
rect 5977 3290 5983 3292
rect 6039 3290 6063 3292
rect 6119 3290 6143 3292
rect 6199 3290 6223 3292
rect 6279 3290 6285 3292
rect 6039 3238 6041 3290
rect 6221 3238 6223 3290
rect 5977 3236 5983 3238
rect 6039 3236 6063 3238
rect 6119 3236 6143 3238
rect 6199 3236 6223 3238
rect 6279 3236 6285 3238
rect 5977 3227 6285 3236
rect 6380 3194 6408 3674
rect 6472 3466 6500 3878
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5184 2650 5212 2926
rect 5317 2748 5625 2757
rect 5317 2746 5323 2748
rect 5379 2746 5403 2748
rect 5459 2746 5483 2748
rect 5539 2746 5563 2748
rect 5619 2746 5625 2748
rect 5379 2694 5381 2746
rect 5561 2694 5563 2746
rect 5317 2692 5323 2694
rect 5379 2692 5403 2694
rect 5459 2692 5483 2694
rect 5539 2692 5563 2694
rect 5619 2692 5625 2694
rect 5317 2683 5625 2692
rect 5736 2650 5764 2994
rect 5814 2952 5870 2961
rect 5814 2887 5870 2896
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5828 2446 5856 2887
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6368 2372 6420 2378
rect 6472 2360 6500 3402
rect 6564 3126 6592 7346
rect 6656 6866 6684 7346
rect 6748 6866 6776 7822
rect 6932 7410 6960 7890
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 6920 7404 6972 7410
rect 6840 7364 6920 7392
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6642 6624 6698 6633
rect 6642 6559 6698 6568
rect 6656 6186 6684 6559
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6644 5772 6696 5778
rect 6748 5760 6776 6802
rect 6840 6322 6868 7364
rect 6920 7346 6972 7352
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7024 7188 7052 7346
rect 7116 7206 7144 7754
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 6932 7160 7052 7188
rect 7104 7200 7156 7206
rect 6932 6984 6960 7160
rect 7104 7142 7156 7148
rect 7064 7100 7372 7109
rect 7064 7098 7070 7100
rect 7126 7098 7150 7100
rect 7206 7098 7230 7100
rect 7286 7098 7310 7100
rect 7366 7098 7372 7100
rect 7126 7046 7128 7098
rect 7308 7046 7310 7098
rect 7064 7044 7070 7046
rect 7126 7044 7150 7046
rect 7206 7044 7230 7046
rect 7286 7044 7310 7046
rect 7366 7044 7372 7046
rect 7064 7035 7372 7044
rect 7484 6984 7512 7346
rect 6932 6956 7052 6984
rect 7024 6633 7052 6956
rect 7116 6956 7512 6984
rect 7010 6624 7066 6633
rect 7010 6559 7066 6568
rect 7116 6390 7144 6956
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7196 6724 7248 6730
rect 7248 6684 7328 6712
rect 7196 6666 7248 6672
rect 7104 6384 7156 6390
rect 7156 6344 7236 6372
rect 7104 6326 7156 6332
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 7104 6248 7156 6254
rect 7010 6216 7066 6225
rect 6828 6180 6880 6186
rect 7066 6196 7104 6202
rect 7066 6190 7156 6196
rect 7066 6174 7144 6190
rect 7010 6151 7066 6160
rect 6828 6122 6880 6128
rect 6696 5732 6776 5760
rect 6644 5714 6696 5720
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6656 2582 6684 5510
rect 6748 4826 6776 5732
rect 6840 5574 6868 6122
rect 7208 6118 7236 6344
rect 7300 6202 7328 6684
rect 7380 6384 7432 6390
rect 7484 6372 7512 6802
rect 7432 6344 7512 6372
rect 7380 6326 7432 6332
rect 7300 6174 7512 6202
rect 7012 6112 7064 6118
rect 6932 6072 7012 6100
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6748 3602 6776 4762
rect 6840 4690 6868 5510
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6840 3126 6868 4014
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 6840 2446 6868 2790
rect 6932 2446 6960 6072
rect 7012 6054 7064 6060
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7064 6012 7372 6021
rect 7064 6010 7070 6012
rect 7126 6010 7150 6012
rect 7206 6010 7230 6012
rect 7286 6010 7310 6012
rect 7366 6010 7372 6012
rect 7126 5958 7128 6010
rect 7308 5958 7310 6010
rect 7064 5956 7070 5958
rect 7126 5956 7150 5958
rect 7206 5956 7230 5958
rect 7286 5956 7310 5958
rect 7366 5956 7372 5958
rect 7064 5947 7372 5956
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7392 5234 7420 5782
rect 7484 5370 7512 6174
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7380 5228 7432 5234
rect 7432 5188 7512 5216
rect 7380 5170 7432 5176
rect 7064 4924 7372 4933
rect 7064 4922 7070 4924
rect 7126 4922 7150 4924
rect 7206 4922 7230 4924
rect 7286 4922 7310 4924
rect 7366 4922 7372 4924
rect 7126 4870 7128 4922
rect 7308 4870 7310 4922
rect 7064 4868 7070 4870
rect 7126 4868 7150 4870
rect 7206 4868 7230 4870
rect 7286 4868 7310 4870
rect 7366 4868 7372 4870
rect 7064 4859 7372 4868
rect 7484 4808 7512 5188
rect 7392 4780 7512 4808
rect 7392 4214 7420 4780
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7484 4282 7512 4626
rect 7576 4282 7604 8434
rect 7668 5302 7696 8894
rect 7724 8732 8032 8741
rect 7724 8730 7730 8732
rect 7786 8730 7810 8732
rect 7866 8730 7890 8732
rect 7946 8730 7970 8732
rect 8026 8730 8032 8732
rect 7786 8678 7788 8730
rect 7968 8678 7970 8730
rect 7724 8676 7730 8678
rect 7786 8676 7810 8678
rect 7866 8676 7890 8678
rect 7946 8676 7970 8678
rect 8026 8676 8032 8678
rect 7724 8667 8032 8676
rect 9048 8634 9076 10548
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 7724 7644 8032 7653
rect 7724 7642 7730 7644
rect 7786 7642 7810 7644
rect 7866 7642 7890 7644
rect 7946 7642 7970 7644
rect 8026 7642 8032 7644
rect 7786 7590 7788 7642
rect 7968 7590 7970 7642
rect 7724 7588 7730 7590
rect 7786 7588 7810 7590
rect 7866 7588 7890 7590
rect 7946 7588 7970 7590
rect 8026 7588 8032 7590
rect 7724 7579 8032 7588
rect 8128 7585 8156 7686
rect 8114 7576 8170 7585
rect 8114 7511 8170 7520
rect 7724 6556 8032 6565
rect 7724 6554 7730 6556
rect 7786 6554 7810 6556
rect 7866 6554 7890 6556
rect 7946 6554 7970 6556
rect 8026 6554 8032 6556
rect 7786 6502 7788 6554
rect 7968 6502 7970 6554
rect 7724 6500 7730 6502
rect 7786 6500 7810 6502
rect 7866 6500 7890 6502
rect 7946 6500 7970 6502
rect 8026 6500 8032 6502
rect 7724 6491 8032 6500
rect 8220 6254 8248 7822
rect 8208 6248 8260 6254
rect 8114 6216 8170 6225
rect 7840 6180 7892 6186
rect 8208 6190 8260 6196
rect 8114 6151 8170 6160
rect 7840 6122 7892 6128
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7760 5846 7788 6054
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7852 5710 7880 6122
rect 8128 5914 8156 6151
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7724 5468 8032 5477
rect 7724 5466 7730 5468
rect 7786 5466 7810 5468
rect 7866 5466 7890 5468
rect 7946 5466 7970 5468
rect 8026 5466 8032 5468
rect 7786 5414 7788 5466
rect 7968 5414 7970 5466
rect 7724 5412 7730 5414
rect 7786 5412 7810 5414
rect 7866 5412 7890 5414
rect 7946 5412 7970 5414
rect 8026 5412 8032 5414
rect 7724 5403 8032 5412
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7392 3924 7420 4150
rect 7668 3942 7696 4966
rect 7724 4380 8032 4389
rect 7724 4378 7730 4380
rect 7786 4378 7810 4380
rect 7866 4378 7890 4380
rect 7946 4378 7970 4380
rect 8026 4378 8032 4380
rect 7786 4326 7788 4378
rect 7968 4326 7970 4378
rect 7724 4324 7730 4326
rect 7786 4324 7810 4326
rect 7866 4324 7890 4326
rect 7946 4324 7970 4326
rect 8026 4324 8032 4326
rect 7724 4315 8032 4324
rect 8128 4185 8156 5170
rect 8220 4214 8248 6190
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8208 4208 8260 4214
rect 8114 4176 8170 4185
rect 7748 4140 7800 4146
rect 8208 4150 8260 4156
rect 8114 4111 8170 4120
rect 7748 4082 7800 4088
rect 7656 3936 7708 3942
rect 7392 3896 7604 3924
rect 7064 3836 7372 3845
rect 7064 3834 7070 3836
rect 7126 3834 7150 3836
rect 7206 3834 7230 3836
rect 7286 3834 7310 3836
rect 7366 3834 7372 3836
rect 7126 3782 7128 3834
rect 7308 3782 7310 3834
rect 7064 3780 7070 3782
rect 7126 3780 7150 3782
rect 7206 3780 7230 3782
rect 7286 3780 7310 3782
rect 7366 3780 7372 3782
rect 7064 3771 7372 3780
rect 7576 3738 7604 3896
rect 7656 3878 7708 3884
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7472 3460 7524 3466
rect 7472 3402 7524 3408
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7116 3058 7144 3334
rect 7484 3194 7512 3402
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7576 3126 7604 3674
rect 7760 3466 7788 4082
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7852 3466 7880 4014
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7724 3292 8032 3301
rect 7724 3290 7730 3292
rect 7786 3290 7810 3292
rect 7866 3290 7890 3292
rect 7946 3290 7970 3292
rect 8026 3290 8032 3292
rect 7786 3238 7788 3290
rect 7968 3238 7970 3290
rect 7724 3236 7730 3238
rect 7786 3236 7810 3238
rect 7866 3236 7890 3238
rect 7946 3236 7970 3238
rect 8026 3236 8032 3238
rect 7724 3227 8032 3236
rect 7564 3120 7616 3126
rect 7564 3062 7616 3068
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7064 2748 7372 2757
rect 7064 2746 7070 2748
rect 7126 2746 7150 2748
rect 7206 2746 7230 2748
rect 7286 2746 7310 2748
rect 7366 2746 7372 2748
rect 7126 2694 7128 2746
rect 7308 2694 7310 2746
rect 7064 2692 7070 2694
rect 7126 2692 7150 2694
rect 7206 2692 7230 2694
rect 7286 2692 7310 2694
rect 7366 2692 7372 2694
rect 7064 2683 7372 2692
rect 7668 2650 7696 2994
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 6420 2332 6500 2360
rect 6368 2314 6420 2320
rect 5448 2304 5500 2310
rect 5092 2264 5448 2292
rect 5448 2246 5500 2252
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 5977 2204 6285 2213
rect 5977 2202 5983 2204
rect 6039 2202 6063 2204
rect 6119 2202 6143 2204
rect 6199 2202 6223 2204
rect 6279 2202 6285 2204
rect 6039 2150 6041 2202
rect 6221 2150 6223 2202
rect 5977 2148 5983 2150
rect 6039 2148 6063 2150
rect 6119 2148 6143 2150
rect 6199 2148 6223 2150
rect 6279 2148 6285 2150
rect 5977 2139 6285 2148
rect 5000 1142 5212 1170
rect 5184 800 5212 1142
rect 6472 870 6592 898
rect 6472 800 6500 870
rect 3330 776 3386 785
rect 3330 711 3386 720
rect 4158 776 4214 785
rect 4158 711 4214 720
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 6564 762 6592 870
rect 6840 762 6868 2246
rect 7724 2204 8032 2213
rect 7724 2202 7730 2204
rect 7786 2202 7810 2204
rect 7866 2202 7890 2204
rect 7946 2202 7970 2204
rect 8026 2202 8032 2204
rect 7786 2150 7788 2202
rect 7968 2150 7970 2202
rect 7724 2148 7730 2150
rect 7786 2148 7810 2150
rect 7866 2148 7890 2150
rect 7946 2148 7970 2150
rect 8026 2148 8032 2150
rect 7724 2139 8032 2148
rect 8404 800 8432 4490
rect 6564 734 6868 762
rect 8390 0 8446 800
<< via2 >>
rect 2778 10240 2834 10296
rect 1490 8880 1546 8936
rect 2489 8730 2545 8732
rect 2569 8730 2625 8732
rect 2649 8730 2705 8732
rect 2729 8730 2785 8732
rect 2489 8678 2535 8730
rect 2535 8678 2545 8730
rect 2569 8678 2599 8730
rect 2599 8678 2611 8730
rect 2611 8678 2625 8730
rect 2649 8678 2663 8730
rect 2663 8678 2675 8730
rect 2675 8678 2705 8730
rect 2729 8678 2739 8730
rect 2739 8678 2785 8730
rect 2489 8676 2545 8678
rect 2569 8676 2625 8678
rect 2649 8676 2705 8678
rect 2729 8676 2785 8678
rect 1829 8186 1885 8188
rect 1909 8186 1965 8188
rect 1989 8186 2045 8188
rect 2069 8186 2125 8188
rect 1829 8134 1875 8186
rect 1875 8134 1885 8186
rect 1909 8134 1939 8186
rect 1939 8134 1951 8186
rect 1951 8134 1965 8186
rect 1989 8134 2003 8186
rect 2003 8134 2015 8186
rect 2015 8134 2045 8186
rect 2069 8134 2079 8186
rect 2079 8134 2125 8186
rect 1829 8132 1885 8134
rect 1909 8132 1965 8134
rect 1989 8132 2045 8134
rect 2069 8132 2125 8134
rect 2686 7828 2688 7848
rect 2688 7828 2740 7848
rect 2740 7828 2742 7848
rect 938 6860 994 6896
rect 938 6840 940 6860
rect 940 6840 992 6860
rect 992 6840 994 6860
rect 1214 6704 1270 6760
rect 938 4800 994 4856
rect 1829 7098 1885 7100
rect 1909 7098 1965 7100
rect 1989 7098 2045 7100
rect 2069 7098 2125 7100
rect 1829 7046 1875 7098
rect 1875 7046 1885 7098
rect 1909 7046 1939 7098
rect 1939 7046 1951 7098
rect 1951 7046 1965 7098
rect 1989 7046 2003 7098
rect 2003 7046 2015 7098
rect 2015 7046 2045 7098
rect 2069 7046 2079 7098
rect 2079 7046 2125 7098
rect 1829 7044 1885 7046
rect 1909 7044 1965 7046
rect 1989 7044 2045 7046
rect 2069 7044 2125 7046
rect 2686 7792 2742 7828
rect 2489 7642 2545 7644
rect 2569 7642 2625 7644
rect 2649 7642 2705 7644
rect 2729 7642 2785 7644
rect 2489 7590 2535 7642
rect 2535 7590 2545 7642
rect 2569 7590 2599 7642
rect 2599 7590 2611 7642
rect 2611 7590 2625 7642
rect 2649 7590 2663 7642
rect 2663 7590 2675 7642
rect 2675 7590 2705 7642
rect 2729 7590 2739 7642
rect 2739 7590 2785 7642
rect 2489 7588 2545 7590
rect 2569 7588 2625 7590
rect 2649 7588 2705 7590
rect 2729 7588 2785 7590
rect 2226 6296 2282 6352
rect 1829 6010 1885 6012
rect 1909 6010 1965 6012
rect 1989 6010 2045 6012
rect 2069 6010 2125 6012
rect 1829 5958 1875 6010
rect 1875 5958 1885 6010
rect 1909 5958 1939 6010
rect 1939 5958 1951 6010
rect 1951 5958 1965 6010
rect 1989 5958 2003 6010
rect 2003 5958 2015 6010
rect 2015 5958 2045 6010
rect 2069 5958 2079 6010
rect 2079 5958 2125 6010
rect 1829 5956 1885 5958
rect 1909 5956 1965 5958
rect 1989 5956 2045 5958
rect 2069 5956 2125 5958
rect 2686 6976 2742 7032
rect 2686 6704 2742 6760
rect 2489 6554 2545 6556
rect 2569 6554 2625 6556
rect 2649 6554 2705 6556
rect 2729 6554 2785 6556
rect 2489 6502 2535 6554
rect 2535 6502 2545 6554
rect 2569 6502 2599 6554
rect 2599 6502 2611 6554
rect 2611 6502 2625 6554
rect 2649 6502 2663 6554
rect 2663 6502 2675 6554
rect 2675 6502 2705 6554
rect 2729 6502 2739 6554
rect 2739 6502 2785 6554
rect 2489 6500 2545 6502
rect 2569 6500 2625 6502
rect 2649 6500 2705 6502
rect 2729 6500 2785 6502
rect 4236 8730 4292 8732
rect 4316 8730 4372 8732
rect 4396 8730 4452 8732
rect 4476 8730 4532 8732
rect 4236 8678 4282 8730
rect 4282 8678 4292 8730
rect 4316 8678 4346 8730
rect 4346 8678 4358 8730
rect 4358 8678 4372 8730
rect 4396 8678 4410 8730
rect 4410 8678 4422 8730
rect 4422 8678 4452 8730
rect 4476 8678 4486 8730
rect 4486 8678 4532 8730
rect 4236 8676 4292 8678
rect 4316 8676 4372 8678
rect 4396 8676 4452 8678
rect 4476 8676 4532 8678
rect 3576 8186 3632 8188
rect 3656 8186 3712 8188
rect 3736 8186 3792 8188
rect 3816 8186 3872 8188
rect 3576 8134 3622 8186
rect 3622 8134 3632 8186
rect 3656 8134 3686 8186
rect 3686 8134 3698 8186
rect 3698 8134 3712 8186
rect 3736 8134 3750 8186
rect 3750 8134 3762 8186
rect 3762 8134 3792 8186
rect 3816 8134 3826 8186
rect 3826 8134 3872 8186
rect 3576 8132 3632 8134
rect 3656 8132 3712 8134
rect 3736 8132 3792 8134
rect 3816 8132 3872 8134
rect 3146 6976 3202 7032
rect 1829 4922 1885 4924
rect 1909 4922 1965 4924
rect 1989 4922 2045 4924
rect 2069 4922 2125 4924
rect 1829 4870 1875 4922
rect 1875 4870 1885 4922
rect 1909 4870 1939 4922
rect 1939 4870 1951 4922
rect 1951 4870 1965 4922
rect 1989 4870 2003 4922
rect 2003 4870 2015 4922
rect 2015 4870 2045 4922
rect 2069 4870 2079 4922
rect 2079 4870 2125 4922
rect 1829 4868 1885 4870
rect 1909 4868 1965 4870
rect 1989 4868 2045 4870
rect 2069 4868 2125 4870
rect 1829 3834 1885 3836
rect 1909 3834 1965 3836
rect 1989 3834 2045 3836
rect 2069 3834 2125 3836
rect 1829 3782 1875 3834
rect 1875 3782 1885 3834
rect 1909 3782 1939 3834
rect 1939 3782 1951 3834
rect 1951 3782 1965 3834
rect 1989 3782 2003 3834
rect 2003 3782 2015 3834
rect 2015 3782 2045 3834
rect 2069 3782 2079 3834
rect 2079 3782 2125 3834
rect 1829 3780 1885 3782
rect 1909 3780 1965 3782
rect 1989 3780 2045 3782
rect 2069 3780 2125 3782
rect 2134 2896 2190 2952
rect 1829 2746 1885 2748
rect 1909 2746 1965 2748
rect 1989 2746 2045 2748
rect 2069 2746 2125 2748
rect 1829 2694 1875 2746
rect 1875 2694 1885 2746
rect 1909 2694 1939 2746
rect 1939 2694 1951 2746
rect 1951 2694 1965 2746
rect 1989 2694 2003 2746
rect 2003 2694 2015 2746
rect 2015 2694 2045 2746
rect 2069 2694 2079 2746
rect 2079 2694 2125 2746
rect 1829 2692 1885 2694
rect 1909 2692 1965 2694
rect 1989 2692 2045 2694
rect 2069 2692 2125 2694
rect 2489 5466 2545 5468
rect 2569 5466 2625 5468
rect 2649 5466 2705 5468
rect 2729 5466 2785 5468
rect 2489 5414 2535 5466
rect 2535 5414 2545 5466
rect 2569 5414 2599 5466
rect 2599 5414 2611 5466
rect 2611 5414 2625 5466
rect 2649 5414 2663 5466
rect 2663 5414 2675 5466
rect 2675 5414 2705 5466
rect 2729 5414 2739 5466
rect 2739 5414 2785 5466
rect 2489 5412 2545 5414
rect 2569 5412 2625 5414
rect 2649 5412 2705 5414
rect 2729 5412 2785 5414
rect 2778 5072 2834 5128
rect 2489 4378 2545 4380
rect 2569 4378 2625 4380
rect 2649 4378 2705 4380
rect 2729 4378 2785 4380
rect 2489 4326 2535 4378
rect 2535 4326 2545 4378
rect 2569 4326 2599 4378
rect 2599 4326 2611 4378
rect 2611 4326 2625 4378
rect 2649 4326 2663 4378
rect 2663 4326 2675 4378
rect 2675 4326 2705 4378
rect 2729 4326 2739 4378
rect 2739 4326 2785 4378
rect 2489 4324 2545 4326
rect 2569 4324 2625 4326
rect 2649 4324 2705 4326
rect 2729 4324 2785 4326
rect 7102 9560 7158 9616
rect 5983 8730 6039 8732
rect 6063 8730 6119 8732
rect 6143 8730 6199 8732
rect 6223 8730 6279 8732
rect 5983 8678 6029 8730
rect 6029 8678 6039 8730
rect 6063 8678 6093 8730
rect 6093 8678 6105 8730
rect 6105 8678 6119 8730
rect 6143 8678 6157 8730
rect 6157 8678 6169 8730
rect 6169 8678 6199 8730
rect 6223 8678 6233 8730
rect 6233 8678 6279 8730
rect 5983 8676 6039 8678
rect 6063 8676 6119 8678
rect 6143 8676 6199 8678
rect 6223 8676 6279 8678
rect 4236 7642 4292 7644
rect 4316 7642 4372 7644
rect 4396 7642 4452 7644
rect 4476 7642 4532 7644
rect 4236 7590 4282 7642
rect 4282 7590 4292 7642
rect 4316 7590 4346 7642
rect 4346 7590 4358 7642
rect 4358 7590 4372 7642
rect 4396 7590 4410 7642
rect 4410 7590 4422 7642
rect 4422 7590 4452 7642
rect 4476 7590 4486 7642
rect 4486 7590 4532 7642
rect 4236 7588 4292 7590
rect 4316 7588 4372 7590
rect 4396 7588 4452 7590
rect 4476 7588 4532 7590
rect 3576 7098 3632 7100
rect 3656 7098 3712 7100
rect 3736 7098 3792 7100
rect 3816 7098 3872 7100
rect 3576 7046 3622 7098
rect 3622 7046 3632 7098
rect 3656 7046 3686 7098
rect 3686 7046 3698 7098
rect 3698 7046 3712 7098
rect 3736 7046 3750 7098
rect 3750 7046 3762 7098
rect 3762 7046 3792 7098
rect 3816 7046 3826 7098
rect 3826 7046 3872 7098
rect 3576 7044 3632 7046
rect 3656 7044 3712 7046
rect 3736 7044 3792 7046
rect 3816 7044 3872 7046
rect 2489 3290 2545 3292
rect 2569 3290 2625 3292
rect 2649 3290 2705 3292
rect 2729 3290 2785 3292
rect 2489 3238 2535 3290
rect 2535 3238 2545 3290
rect 2569 3238 2599 3290
rect 2599 3238 2611 3290
rect 2611 3238 2625 3290
rect 2649 3238 2663 3290
rect 2663 3238 2675 3290
rect 2675 3238 2705 3290
rect 2729 3238 2739 3290
rect 2739 3238 2785 3290
rect 2489 3236 2545 3238
rect 2569 3236 2625 3238
rect 2649 3236 2705 3238
rect 2729 3236 2785 3238
rect 3576 6010 3632 6012
rect 3656 6010 3712 6012
rect 3736 6010 3792 6012
rect 3816 6010 3872 6012
rect 3576 5958 3622 6010
rect 3622 5958 3632 6010
rect 3656 5958 3686 6010
rect 3686 5958 3698 6010
rect 3698 5958 3712 6010
rect 3736 5958 3750 6010
rect 3750 5958 3762 6010
rect 3762 5958 3792 6010
rect 3816 5958 3826 6010
rect 3826 5958 3872 6010
rect 3576 5956 3632 5958
rect 3656 5956 3712 5958
rect 3736 5956 3792 5958
rect 3816 5956 3872 5958
rect 4236 6554 4292 6556
rect 4316 6554 4372 6556
rect 4396 6554 4452 6556
rect 4476 6554 4532 6556
rect 4236 6502 4282 6554
rect 4282 6502 4292 6554
rect 4316 6502 4346 6554
rect 4346 6502 4358 6554
rect 4358 6502 4372 6554
rect 4396 6502 4410 6554
rect 4410 6502 4422 6554
rect 4422 6502 4452 6554
rect 4476 6502 4486 6554
rect 4486 6502 4532 6554
rect 4236 6500 4292 6502
rect 4316 6500 4372 6502
rect 4396 6500 4452 6502
rect 4476 6500 4532 6502
rect 3576 4922 3632 4924
rect 3656 4922 3712 4924
rect 3736 4922 3792 4924
rect 3816 4922 3872 4924
rect 3576 4870 3622 4922
rect 3622 4870 3632 4922
rect 3656 4870 3686 4922
rect 3686 4870 3698 4922
rect 3698 4870 3712 4922
rect 3736 4870 3750 4922
rect 3750 4870 3762 4922
rect 3762 4870 3792 4922
rect 3816 4870 3826 4922
rect 3826 4870 3872 4922
rect 3576 4868 3632 4870
rect 3656 4868 3712 4870
rect 3736 4868 3792 4870
rect 3816 4868 3872 4870
rect 3514 3984 3570 4040
rect 3576 3834 3632 3836
rect 3656 3834 3712 3836
rect 3736 3834 3792 3836
rect 3816 3834 3872 3836
rect 3576 3782 3622 3834
rect 3622 3782 3632 3834
rect 3656 3782 3686 3834
rect 3686 3782 3698 3834
rect 3698 3782 3712 3834
rect 3736 3782 3750 3834
rect 3750 3782 3762 3834
rect 3762 3782 3792 3834
rect 3816 3782 3826 3834
rect 3826 3782 3872 3834
rect 3576 3780 3632 3782
rect 3656 3780 3712 3782
rect 3736 3780 3792 3782
rect 3816 3780 3872 3782
rect 4236 5466 4292 5468
rect 4316 5466 4372 5468
rect 4396 5466 4452 5468
rect 4476 5466 4532 5468
rect 4236 5414 4282 5466
rect 4282 5414 4292 5466
rect 4316 5414 4346 5466
rect 4346 5414 4358 5466
rect 4358 5414 4372 5466
rect 4396 5414 4410 5466
rect 4410 5414 4422 5466
rect 4422 5414 4452 5466
rect 4476 5414 4486 5466
rect 4486 5414 4532 5466
rect 4236 5412 4292 5414
rect 4316 5412 4372 5414
rect 4396 5412 4452 5414
rect 4476 5412 4532 5414
rect 2489 2202 2545 2204
rect 2569 2202 2625 2204
rect 2649 2202 2705 2204
rect 2729 2202 2785 2204
rect 2489 2150 2535 2202
rect 2535 2150 2545 2202
rect 2569 2150 2599 2202
rect 2599 2150 2611 2202
rect 2611 2150 2625 2202
rect 2649 2150 2663 2202
rect 2663 2150 2675 2202
rect 2675 2150 2705 2202
rect 2729 2150 2739 2202
rect 2739 2150 2785 2202
rect 2489 2148 2545 2150
rect 2569 2148 2625 2150
rect 2649 2148 2705 2150
rect 2729 2148 2785 2150
rect 3576 2746 3632 2748
rect 3656 2746 3712 2748
rect 3736 2746 3792 2748
rect 3816 2746 3872 2748
rect 3576 2694 3622 2746
rect 3622 2694 3632 2746
rect 3656 2694 3686 2746
rect 3686 2694 3698 2746
rect 3698 2694 3712 2746
rect 3736 2694 3750 2746
rect 3750 2694 3762 2746
rect 3762 2694 3792 2746
rect 3816 2694 3826 2746
rect 3826 2694 3872 2746
rect 3576 2692 3632 2694
rect 3656 2692 3712 2694
rect 3736 2692 3792 2694
rect 3816 2692 3872 2694
rect 4236 4378 4292 4380
rect 4316 4378 4372 4380
rect 4396 4378 4452 4380
rect 4476 4378 4532 4380
rect 4236 4326 4282 4378
rect 4282 4326 4292 4378
rect 4316 4326 4346 4378
rect 4346 4326 4358 4378
rect 4358 4326 4372 4378
rect 4396 4326 4410 4378
rect 4410 4326 4422 4378
rect 4422 4326 4452 4378
rect 4476 4326 4486 4378
rect 4486 4326 4532 4378
rect 4236 4324 4292 4326
rect 4316 4324 4372 4326
rect 4396 4324 4452 4326
rect 4476 4324 4532 4326
rect 4236 3290 4292 3292
rect 4316 3290 4372 3292
rect 4396 3290 4452 3292
rect 4476 3290 4532 3292
rect 4236 3238 4282 3290
rect 4282 3238 4292 3290
rect 4316 3238 4346 3290
rect 4346 3238 4358 3290
rect 4358 3238 4372 3290
rect 4396 3238 4410 3290
rect 4410 3238 4422 3290
rect 4422 3238 4452 3290
rect 4476 3238 4486 3290
rect 4486 3238 4532 3290
rect 4236 3236 4292 3238
rect 4316 3236 4372 3238
rect 4396 3236 4452 3238
rect 4476 3236 4532 3238
rect 3146 1400 3202 1456
rect 5323 8186 5379 8188
rect 5403 8186 5459 8188
rect 5483 8186 5539 8188
rect 5563 8186 5619 8188
rect 5323 8134 5369 8186
rect 5369 8134 5379 8186
rect 5403 8134 5433 8186
rect 5433 8134 5445 8186
rect 5445 8134 5459 8186
rect 5483 8134 5497 8186
rect 5497 8134 5509 8186
rect 5509 8134 5539 8186
rect 5563 8134 5573 8186
rect 5573 8134 5619 8186
rect 5323 8132 5379 8134
rect 5403 8132 5459 8134
rect 5483 8132 5539 8134
rect 5563 8132 5619 8134
rect 5262 7792 5318 7848
rect 5983 7642 6039 7644
rect 6063 7642 6119 7644
rect 6143 7642 6199 7644
rect 6223 7642 6279 7644
rect 5983 7590 6029 7642
rect 6029 7590 6039 7642
rect 6063 7590 6093 7642
rect 6093 7590 6105 7642
rect 6105 7590 6119 7642
rect 6143 7590 6157 7642
rect 6157 7590 6169 7642
rect 6169 7590 6199 7642
rect 6223 7590 6233 7642
rect 6233 7590 6279 7642
rect 5983 7588 6039 7590
rect 6063 7588 6119 7590
rect 6143 7588 6199 7590
rect 6223 7588 6279 7590
rect 7070 8186 7126 8188
rect 7150 8186 7206 8188
rect 7230 8186 7286 8188
rect 7310 8186 7366 8188
rect 7070 8134 7116 8186
rect 7116 8134 7126 8186
rect 7150 8134 7180 8186
rect 7180 8134 7192 8186
rect 7192 8134 7206 8186
rect 7230 8134 7244 8186
rect 7244 8134 7256 8186
rect 7256 8134 7286 8186
rect 7310 8134 7320 8186
rect 7320 8134 7366 8186
rect 7070 8132 7126 8134
rect 7150 8132 7206 8134
rect 7230 8132 7286 8134
rect 7310 8132 7366 8134
rect 5323 7098 5379 7100
rect 5403 7098 5459 7100
rect 5483 7098 5539 7100
rect 5563 7098 5619 7100
rect 5323 7046 5369 7098
rect 5369 7046 5379 7098
rect 5403 7046 5433 7098
rect 5433 7046 5445 7098
rect 5445 7046 5459 7098
rect 5483 7046 5497 7098
rect 5497 7046 5509 7098
rect 5509 7046 5539 7098
rect 5563 7046 5573 7098
rect 5573 7046 5619 7098
rect 5323 7044 5379 7046
rect 5403 7044 5459 7046
rect 5483 7044 5539 7046
rect 5563 7044 5619 7046
rect 5323 6010 5379 6012
rect 5403 6010 5459 6012
rect 5483 6010 5539 6012
rect 5563 6010 5619 6012
rect 5323 5958 5369 6010
rect 5369 5958 5379 6010
rect 5403 5958 5433 6010
rect 5433 5958 5445 6010
rect 5445 5958 5459 6010
rect 5483 5958 5497 6010
rect 5497 5958 5509 6010
rect 5509 5958 5539 6010
rect 5563 5958 5573 6010
rect 5573 5958 5619 6010
rect 5323 5956 5379 5958
rect 5403 5956 5459 5958
rect 5483 5956 5539 5958
rect 5563 5956 5619 5958
rect 5323 4922 5379 4924
rect 5403 4922 5459 4924
rect 5483 4922 5539 4924
rect 5563 4922 5619 4924
rect 5323 4870 5369 4922
rect 5369 4870 5379 4922
rect 5403 4870 5433 4922
rect 5433 4870 5445 4922
rect 5445 4870 5459 4922
rect 5483 4870 5497 4922
rect 5497 4870 5509 4922
rect 5509 4870 5539 4922
rect 5563 4870 5573 4922
rect 5573 4870 5619 4922
rect 5323 4868 5379 4870
rect 5403 4868 5459 4870
rect 5483 4868 5539 4870
rect 5563 4868 5619 4870
rect 5983 6554 6039 6556
rect 6063 6554 6119 6556
rect 6143 6554 6199 6556
rect 6223 6554 6279 6556
rect 5983 6502 6029 6554
rect 6029 6502 6039 6554
rect 6063 6502 6093 6554
rect 6093 6502 6105 6554
rect 6105 6502 6119 6554
rect 6143 6502 6157 6554
rect 6157 6502 6169 6554
rect 6169 6502 6199 6554
rect 6223 6502 6233 6554
rect 6233 6502 6279 6554
rect 5983 6500 6039 6502
rect 6063 6500 6119 6502
rect 6143 6500 6199 6502
rect 6223 6500 6279 6502
rect 6366 6160 6422 6216
rect 5983 5466 6039 5468
rect 6063 5466 6119 5468
rect 6143 5466 6199 5468
rect 6223 5466 6279 5468
rect 5983 5414 6029 5466
rect 6029 5414 6039 5466
rect 6063 5414 6093 5466
rect 6093 5414 6105 5466
rect 6105 5414 6119 5466
rect 6143 5414 6157 5466
rect 6157 5414 6169 5466
rect 6169 5414 6199 5466
rect 6223 5414 6233 5466
rect 6233 5414 6279 5466
rect 5983 5412 6039 5414
rect 6063 5412 6119 5414
rect 6143 5412 6199 5414
rect 6223 5412 6279 5414
rect 4236 2202 4292 2204
rect 4316 2202 4372 2204
rect 4396 2202 4452 2204
rect 4476 2202 4532 2204
rect 4236 2150 4282 2202
rect 4282 2150 4292 2202
rect 4316 2150 4346 2202
rect 4346 2150 4358 2202
rect 4358 2150 4372 2202
rect 4396 2150 4410 2202
rect 4410 2150 4422 2202
rect 4422 2150 4452 2202
rect 4476 2150 4486 2202
rect 4486 2150 4532 2202
rect 4236 2148 4292 2150
rect 4316 2148 4372 2150
rect 4396 2148 4452 2150
rect 4476 2148 4532 2150
rect 4894 2352 4950 2408
rect 5323 3834 5379 3836
rect 5403 3834 5459 3836
rect 5483 3834 5539 3836
rect 5563 3834 5619 3836
rect 5323 3782 5369 3834
rect 5369 3782 5379 3834
rect 5403 3782 5433 3834
rect 5433 3782 5445 3834
rect 5445 3782 5459 3834
rect 5483 3782 5497 3834
rect 5497 3782 5509 3834
rect 5509 3782 5539 3834
rect 5563 3782 5573 3834
rect 5573 3782 5619 3834
rect 5323 3780 5379 3782
rect 5403 3780 5459 3782
rect 5483 3780 5539 3782
rect 5563 3780 5619 3782
rect 5983 4378 6039 4380
rect 6063 4378 6119 4380
rect 6143 4378 6199 4380
rect 6223 4378 6279 4380
rect 5983 4326 6029 4378
rect 6029 4326 6039 4378
rect 6063 4326 6093 4378
rect 6093 4326 6105 4378
rect 6105 4326 6119 4378
rect 6143 4326 6157 4378
rect 6157 4326 6169 4378
rect 6169 4326 6199 4378
rect 6223 4326 6233 4378
rect 6233 4326 6279 4378
rect 5983 4324 6039 4326
rect 6063 4324 6119 4326
rect 6143 4324 6199 4326
rect 6223 4324 6279 4326
rect 5983 3290 6039 3292
rect 6063 3290 6119 3292
rect 6143 3290 6199 3292
rect 6223 3290 6279 3292
rect 5983 3238 6029 3290
rect 6029 3238 6039 3290
rect 6063 3238 6093 3290
rect 6093 3238 6105 3290
rect 6105 3238 6119 3290
rect 6143 3238 6157 3290
rect 6157 3238 6169 3290
rect 6169 3238 6199 3290
rect 6223 3238 6233 3290
rect 6233 3238 6279 3290
rect 5983 3236 6039 3238
rect 6063 3236 6119 3238
rect 6143 3236 6199 3238
rect 6223 3236 6279 3238
rect 5323 2746 5379 2748
rect 5403 2746 5459 2748
rect 5483 2746 5539 2748
rect 5563 2746 5619 2748
rect 5323 2694 5369 2746
rect 5369 2694 5379 2746
rect 5403 2694 5433 2746
rect 5433 2694 5445 2746
rect 5445 2694 5459 2746
rect 5483 2694 5497 2746
rect 5497 2694 5509 2746
rect 5509 2694 5539 2746
rect 5563 2694 5573 2746
rect 5573 2694 5619 2746
rect 5323 2692 5379 2694
rect 5403 2692 5459 2694
rect 5483 2692 5539 2694
rect 5563 2692 5619 2694
rect 5814 2896 5870 2952
rect 6642 6568 6698 6624
rect 7070 7098 7126 7100
rect 7150 7098 7206 7100
rect 7230 7098 7286 7100
rect 7310 7098 7366 7100
rect 7070 7046 7116 7098
rect 7116 7046 7126 7098
rect 7150 7046 7180 7098
rect 7180 7046 7192 7098
rect 7192 7046 7206 7098
rect 7230 7046 7244 7098
rect 7244 7046 7256 7098
rect 7256 7046 7286 7098
rect 7310 7046 7320 7098
rect 7320 7046 7366 7098
rect 7070 7044 7126 7046
rect 7150 7044 7206 7046
rect 7230 7044 7286 7046
rect 7310 7044 7366 7046
rect 7010 6568 7066 6624
rect 7010 6160 7066 6216
rect 7070 6010 7126 6012
rect 7150 6010 7206 6012
rect 7230 6010 7286 6012
rect 7310 6010 7366 6012
rect 7070 5958 7116 6010
rect 7116 5958 7126 6010
rect 7150 5958 7180 6010
rect 7180 5958 7192 6010
rect 7192 5958 7206 6010
rect 7230 5958 7244 6010
rect 7244 5958 7256 6010
rect 7256 5958 7286 6010
rect 7310 5958 7320 6010
rect 7320 5958 7366 6010
rect 7070 5956 7126 5958
rect 7150 5956 7206 5958
rect 7230 5956 7286 5958
rect 7310 5956 7366 5958
rect 7070 4922 7126 4924
rect 7150 4922 7206 4924
rect 7230 4922 7286 4924
rect 7310 4922 7366 4924
rect 7070 4870 7116 4922
rect 7116 4870 7126 4922
rect 7150 4870 7180 4922
rect 7180 4870 7192 4922
rect 7192 4870 7206 4922
rect 7230 4870 7244 4922
rect 7244 4870 7256 4922
rect 7256 4870 7286 4922
rect 7310 4870 7320 4922
rect 7320 4870 7366 4922
rect 7070 4868 7126 4870
rect 7150 4868 7206 4870
rect 7230 4868 7286 4870
rect 7310 4868 7366 4870
rect 7730 8730 7786 8732
rect 7810 8730 7866 8732
rect 7890 8730 7946 8732
rect 7970 8730 8026 8732
rect 7730 8678 7776 8730
rect 7776 8678 7786 8730
rect 7810 8678 7840 8730
rect 7840 8678 7852 8730
rect 7852 8678 7866 8730
rect 7890 8678 7904 8730
rect 7904 8678 7916 8730
rect 7916 8678 7946 8730
rect 7970 8678 7980 8730
rect 7980 8678 8026 8730
rect 7730 8676 7786 8678
rect 7810 8676 7866 8678
rect 7890 8676 7946 8678
rect 7970 8676 8026 8678
rect 7730 7642 7786 7644
rect 7810 7642 7866 7644
rect 7890 7642 7946 7644
rect 7970 7642 8026 7644
rect 7730 7590 7776 7642
rect 7776 7590 7786 7642
rect 7810 7590 7840 7642
rect 7840 7590 7852 7642
rect 7852 7590 7866 7642
rect 7890 7590 7904 7642
rect 7904 7590 7916 7642
rect 7916 7590 7946 7642
rect 7970 7590 7980 7642
rect 7980 7590 8026 7642
rect 7730 7588 7786 7590
rect 7810 7588 7866 7590
rect 7890 7588 7946 7590
rect 7970 7588 8026 7590
rect 8114 7520 8170 7576
rect 7730 6554 7786 6556
rect 7810 6554 7866 6556
rect 7890 6554 7946 6556
rect 7970 6554 8026 6556
rect 7730 6502 7776 6554
rect 7776 6502 7786 6554
rect 7810 6502 7840 6554
rect 7840 6502 7852 6554
rect 7852 6502 7866 6554
rect 7890 6502 7904 6554
rect 7904 6502 7916 6554
rect 7916 6502 7946 6554
rect 7970 6502 7980 6554
rect 7980 6502 8026 6554
rect 7730 6500 7786 6502
rect 7810 6500 7866 6502
rect 7890 6500 7946 6502
rect 7970 6500 8026 6502
rect 8114 6160 8170 6216
rect 7730 5466 7786 5468
rect 7810 5466 7866 5468
rect 7890 5466 7946 5468
rect 7970 5466 8026 5468
rect 7730 5414 7776 5466
rect 7776 5414 7786 5466
rect 7810 5414 7840 5466
rect 7840 5414 7852 5466
rect 7852 5414 7866 5466
rect 7890 5414 7904 5466
rect 7904 5414 7916 5466
rect 7916 5414 7946 5466
rect 7970 5414 7980 5466
rect 7980 5414 8026 5466
rect 7730 5412 7786 5414
rect 7810 5412 7866 5414
rect 7890 5412 7946 5414
rect 7970 5412 8026 5414
rect 7730 4378 7786 4380
rect 7810 4378 7866 4380
rect 7890 4378 7946 4380
rect 7970 4378 8026 4380
rect 7730 4326 7776 4378
rect 7776 4326 7786 4378
rect 7810 4326 7840 4378
rect 7840 4326 7852 4378
rect 7852 4326 7866 4378
rect 7890 4326 7904 4378
rect 7904 4326 7916 4378
rect 7916 4326 7946 4378
rect 7970 4326 7980 4378
rect 7980 4326 8026 4378
rect 7730 4324 7786 4326
rect 7810 4324 7866 4326
rect 7890 4324 7946 4326
rect 7970 4324 8026 4326
rect 8114 4120 8170 4176
rect 7070 3834 7126 3836
rect 7150 3834 7206 3836
rect 7230 3834 7286 3836
rect 7310 3834 7366 3836
rect 7070 3782 7116 3834
rect 7116 3782 7126 3834
rect 7150 3782 7180 3834
rect 7180 3782 7192 3834
rect 7192 3782 7206 3834
rect 7230 3782 7244 3834
rect 7244 3782 7256 3834
rect 7256 3782 7286 3834
rect 7310 3782 7320 3834
rect 7320 3782 7366 3834
rect 7070 3780 7126 3782
rect 7150 3780 7206 3782
rect 7230 3780 7286 3782
rect 7310 3780 7366 3782
rect 7730 3290 7786 3292
rect 7810 3290 7866 3292
rect 7890 3290 7946 3292
rect 7970 3290 8026 3292
rect 7730 3238 7776 3290
rect 7776 3238 7786 3290
rect 7810 3238 7840 3290
rect 7840 3238 7852 3290
rect 7852 3238 7866 3290
rect 7890 3238 7904 3290
rect 7904 3238 7916 3290
rect 7916 3238 7946 3290
rect 7970 3238 7980 3290
rect 7980 3238 8026 3290
rect 7730 3236 7786 3238
rect 7810 3236 7866 3238
rect 7890 3236 7946 3238
rect 7970 3236 8026 3238
rect 7070 2746 7126 2748
rect 7150 2746 7206 2748
rect 7230 2746 7286 2748
rect 7310 2746 7366 2748
rect 7070 2694 7116 2746
rect 7116 2694 7126 2746
rect 7150 2694 7180 2746
rect 7180 2694 7192 2746
rect 7192 2694 7206 2746
rect 7230 2694 7244 2746
rect 7244 2694 7256 2746
rect 7256 2694 7286 2746
rect 7310 2694 7320 2746
rect 7320 2694 7366 2746
rect 7070 2692 7126 2694
rect 7150 2692 7206 2694
rect 7230 2692 7286 2694
rect 7310 2692 7366 2694
rect 5983 2202 6039 2204
rect 6063 2202 6119 2204
rect 6143 2202 6199 2204
rect 6223 2202 6279 2204
rect 5983 2150 6029 2202
rect 6029 2150 6039 2202
rect 6063 2150 6093 2202
rect 6093 2150 6105 2202
rect 6105 2150 6119 2202
rect 6143 2150 6157 2202
rect 6157 2150 6169 2202
rect 6169 2150 6199 2202
rect 6223 2150 6233 2202
rect 6233 2150 6279 2202
rect 5983 2148 6039 2150
rect 6063 2148 6119 2150
rect 6143 2148 6199 2150
rect 6223 2148 6279 2150
rect 3330 720 3386 776
rect 4158 720 4214 776
rect 7730 2202 7786 2204
rect 7810 2202 7866 2204
rect 7890 2202 7946 2204
rect 7970 2202 8026 2204
rect 7730 2150 7776 2202
rect 7776 2150 7786 2202
rect 7810 2150 7840 2202
rect 7840 2150 7852 2202
rect 7852 2150 7866 2202
rect 7890 2150 7904 2202
rect 7904 2150 7916 2202
rect 7916 2150 7946 2202
rect 7970 2150 7980 2202
rect 7980 2150 8026 2202
rect 7730 2148 7786 2150
rect 7810 2148 7866 2150
rect 7890 2148 7946 2150
rect 7970 2148 8026 2150
<< metal3 >>
rect 0 10298 800 10328
rect 2773 10298 2839 10301
rect 0 10296 2839 10298
rect 0 10240 2778 10296
rect 2834 10240 2839 10296
rect 0 10238 2839 10240
rect 0 10208 800 10238
rect 2773 10235 2839 10238
rect 7097 9618 7163 9621
rect 8404 9618 9204 9648
rect 7097 9616 9204 9618
rect 7097 9560 7102 9616
rect 7158 9560 9204 9616
rect 7097 9558 9204 9560
rect 7097 9555 7163 9558
rect 8404 9528 9204 9558
rect 0 8938 800 8968
rect 1485 8938 1551 8941
rect 0 8936 1551 8938
rect 0 8880 1490 8936
rect 1546 8880 1551 8936
rect 0 8878 1551 8880
rect 0 8848 800 8878
rect 1485 8875 1551 8878
rect 2479 8736 2795 8737
rect 2479 8672 2485 8736
rect 2549 8672 2565 8736
rect 2629 8672 2645 8736
rect 2709 8672 2725 8736
rect 2789 8672 2795 8736
rect 2479 8671 2795 8672
rect 4226 8736 4542 8737
rect 4226 8672 4232 8736
rect 4296 8672 4312 8736
rect 4376 8672 4392 8736
rect 4456 8672 4472 8736
rect 4536 8672 4542 8736
rect 4226 8671 4542 8672
rect 5973 8736 6289 8737
rect 5973 8672 5979 8736
rect 6043 8672 6059 8736
rect 6123 8672 6139 8736
rect 6203 8672 6219 8736
rect 6283 8672 6289 8736
rect 5973 8671 6289 8672
rect 7720 8736 8036 8737
rect 7720 8672 7726 8736
rect 7790 8672 7806 8736
rect 7870 8672 7886 8736
rect 7950 8672 7966 8736
rect 8030 8672 8036 8736
rect 7720 8671 8036 8672
rect 1819 8192 2135 8193
rect 1819 8128 1825 8192
rect 1889 8128 1905 8192
rect 1969 8128 1985 8192
rect 2049 8128 2065 8192
rect 2129 8128 2135 8192
rect 1819 8127 2135 8128
rect 3566 8192 3882 8193
rect 3566 8128 3572 8192
rect 3636 8128 3652 8192
rect 3716 8128 3732 8192
rect 3796 8128 3812 8192
rect 3876 8128 3882 8192
rect 3566 8127 3882 8128
rect 5313 8192 5629 8193
rect 5313 8128 5319 8192
rect 5383 8128 5399 8192
rect 5463 8128 5479 8192
rect 5543 8128 5559 8192
rect 5623 8128 5629 8192
rect 5313 8127 5629 8128
rect 7060 8192 7376 8193
rect 7060 8128 7066 8192
rect 7130 8128 7146 8192
rect 7210 8128 7226 8192
rect 7290 8128 7306 8192
rect 7370 8128 7376 8192
rect 7060 8127 7376 8128
rect 2681 7850 2747 7853
rect 5257 7850 5323 7853
rect 2681 7848 5323 7850
rect 2681 7792 2686 7848
rect 2742 7792 5262 7848
rect 5318 7792 5323 7848
rect 2681 7790 5323 7792
rect 2681 7787 2747 7790
rect 5257 7787 5323 7790
rect 2479 7648 2795 7649
rect 2479 7584 2485 7648
rect 2549 7584 2565 7648
rect 2629 7584 2645 7648
rect 2709 7584 2725 7648
rect 2789 7584 2795 7648
rect 2479 7583 2795 7584
rect 4226 7648 4542 7649
rect 4226 7584 4232 7648
rect 4296 7584 4312 7648
rect 4376 7584 4392 7648
rect 4456 7584 4472 7648
rect 4536 7584 4542 7648
rect 4226 7583 4542 7584
rect 5973 7648 6289 7649
rect 5973 7584 5979 7648
rect 6043 7584 6059 7648
rect 6123 7584 6139 7648
rect 6203 7584 6219 7648
rect 6283 7584 6289 7648
rect 5973 7583 6289 7584
rect 7720 7648 8036 7649
rect 7720 7584 7726 7648
rect 7790 7584 7806 7648
rect 7870 7584 7886 7648
rect 7950 7584 7966 7648
rect 8030 7584 8036 7648
rect 7720 7583 8036 7584
rect 8109 7578 8175 7581
rect 8404 7578 9204 7608
rect 8109 7576 9204 7578
rect 8109 7520 8114 7576
rect 8170 7520 9204 7576
rect 8109 7518 9204 7520
rect 8109 7515 8175 7518
rect 8404 7488 9204 7518
rect 1819 7104 2135 7105
rect 1819 7040 1825 7104
rect 1889 7040 1905 7104
rect 1969 7040 1985 7104
rect 2049 7040 2065 7104
rect 2129 7040 2135 7104
rect 1819 7039 2135 7040
rect 3566 7104 3882 7105
rect 3566 7040 3572 7104
rect 3636 7040 3652 7104
rect 3716 7040 3732 7104
rect 3796 7040 3812 7104
rect 3876 7040 3882 7104
rect 3566 7039 3882 7040
rect 5313 7104 5629 7105
rect 5313 7040 5319 7104
rect 5383 7040 5399 7104
rect 5463 7040 5479 7104
rect 5543 7040 5559 7104
rect 5623 7040 5629 7104
rect 5313 7039 5629 7040
rect 7060 7104 7376 7105
rect 7060 7040 7066 7104
rect 7130 7040 7146 7104
rect 7210 7040 7226 7104
rect 7290 7040 7306 7104
rect 7370 7040 7376 7104
rect 7060 7039 7376 7040
rect 2681 7034 2747 7037
rect 3141 7034 3207 7037
rect 2681 7032 3207 7034
rect 2681 6976 2686 7032
rect 2742 6976 3146 7032
rect 3202 6976 3207 7032
rect 2681 6974 3207 6976
rect 2681 6971 2747 6974
rect 3141 6971 3207 6974
rect 0 6898 800 6928
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6808 800 6838
rect 933 6835 999 6838
rect 1209 6762 1275 6765
rect 2681 6762 2747 6765
rect 1209 6760 2747 6762
rect 1209 6704 1214 6760
rect 1270 6704 2686 6760
rect 2742 6704 2747 6760
rect 1209 6702 2747 6704
rect 1209 6699 1275 6702
rect 2681 6699 2747 6702
rect 6637 6626 6703 6629
rect 7005 6626 7071 6629
rect 6637 6624 7071 6626
rect 6637 6568 6642 6624
rect 6698 6568 7010 6624
rect 7066 6568 7071 6624
rect 6637 6566 7071 6568
rect 6637 6563 6703 6566
rect 7005 6563 7071 6566
rect 2479 6560 2795 6561
rect 2479 6496 2485 6560
rect 2549 6496 2565 6560
rect 2629 6496 2645 6560
rect 2709 6496 2725 6560
rect 2789 6496 2795 6560
rect 2479 6495 2795 6496
rect 4226 6560 4542 6561
rect 4226 6496 4232 6560
rect 4296 6496 4312 6560
rect 4376 6496 4392 6560
rect 4456 6496 4472 6560
rect 4536 6496 4542 6560
rect 4226 6495 4542 6496
rect 5973 6560 6289 6561
rect 5973 6496 5979 6560
rect 6043 6496 6059 6560
rect 6123 6496 6139 6560
rect 6203 6496 6219 6560
rect 6283 6496 6289 6560
rect 5973 6495 6289 6496
rect 7720 6560 8036 6561
rect 7720 6496 7726 6560
rect 7790 6496 7806 6560
rect 7870 6496 7886 6560
rect 7950 6496 7966 6560
rect 8030 6496 8036 6560
rect 7720 6495 8036 6496
rect 2221 6356 2287 6357
rect 2221 6352 2268 6356
rect 2332 6354 2338 6356
rect 2221 6296 2226 6352
rect 2221 6292 2268 6296
rect 2332 6294 2378 6354
rect 2332 6292 2338 6294
rect 2221 6291 2287 6292
rect 6361 6218 6427 6221
rect 7005 6218 7071 6221
rect 6361 6216 7071 6218
rect 6361 6160 6366 6216
rect 6422 6160 7010 6216
rect 7066 6160 7071 6216
rect 6361 6158 7071 6160
rect 6361 6155 6427 6158
rect 7005 6155 7071 6158
rect 8109 6218 8175 6221
rect 8404 6218 9204 6248
rect 8109 6216 9204 6218
rect 8109 6160 8114 6216
rect 8170 6160 9204 6216
rect 8109 6158 9204 6160
rect 8109 6155 8175 6158
rect 8404 6128 9204 6158
rect 1819 6016 2135 6017
rect 1819 5952 1825 6016
rect 1889 5952 1905 6016
rect 1969 5952 1985 6016
rect 2049 5952 2065 6016
rect 2129 5952 2135 6016
rect 1819 5951 2135 5952
rect 3566 6016 3882 6017
rect 3566 5952 3572 6016
rect 3636 5952 3652 6016
rect 3716 5952 3732 6016
rect 3796 5952 3812 6016
rect 3876 5952 3882 6016
rect 3566 5951 3882 5952
rect 5313 6016 5629 6017
rect 5313 5952 5319 6016
rect 5383 5952 5399 6016
rect 5463 5952 5479 6016
rect 5543 5952 5559 6016
rect 5623 5952 5629 6016
rect 5313 5951 5629 5952
rect 7060 6016 7376 6017
rect 7060 5952 7066 6016
rect 7130 5952 7146 6016
rect 7210 5952 7226 6016
rect 7290 5952 7306 6016
rect 7370 5952 7376 6016
rect 7060 5951 7376 5952
rect 2479 5472 2795 5473
rect 2479 5408 2485 5472
rect 2549 5408 2565 5472
rect 2629 5408 2645 5472
rect 2709 5408 2725 5472
rect 2789 5408 2795 5472
rect 2479 5407 2795 5408
rect 4226 5472 4542 5473
rect 4226 5408 4232 5472
rect 4296 5408 4312 5472
rect 4376 5408 4392 5472
rect 4456 5408 4472 5472
rect 4536 5408 4542 5472
rect 4226 5407 4542 5408
rect 5973 5472 6289 5473
rect 5973 5408 5979 5472
rect 6043 5408 6059 5472
rect 6123 5408 6139 5472
rect 6203 5408 6219 5472
rect 6283 5408 6289 5472
rect 5973 5407 6289 5408
rect 7720 5472 8036 5473
rect 7720 5408 7726 5472
rect 7790 5408 7806 5472
rect 7870 5408 7886 5472
rect 7950 5408 7966 5472
rect 8030 5408 8036 5472
rect 7720 5407 8036 5408
rect 2773 5130 2839 5133
rect 2998 5130 3004 5132
rect 2773 5128 3004 5130
rect 2773 5072 2778 5128
rect 2834 5072 3004 5128
rect 2773 5070 3004 5072
rect 2773 5067 2839 5070
rect 2998 5068 3004 5070
rect 3068 5068 3074 5132
rect 1819 4928 2135 4929
rect 0 4858 800 4888
rect 1819 4864 1825 4928
rect 1889 4864 1905 4928
rect 1969 4864 1985 4928
rect 2049 4864 2065 4928
rect 2129 4864 2135 4928
rect 1819 4863 2135 4864
rect 3566 4928 3882 4929
rect 3566 4864 3572 4928
rect 3636 4864 3652 4928
rect 3716 4864 3732 4928
rect 3796 4864 3812 4928
rect 3876 4864 3882 4928
rect 3566 4863 3882 4864
rect 5313 4928 5629 4929
rect 5313 4864 5319 4928
rect 5383 4864 5399 4928
rect 5463 4864 5479 4928
rect 5543 4864 5559 4928
rect 5623 4864 5629 4928
rect 5313 4863 5629 4864
rect 7060 4928 7376 4929
rect 7060 4864 7066 4928
rect 7130 4864 7146 4928
rect 7210 4864 7226 4928
rect 7290 4864 7306 4928
rect 7370 4864 7376 4928
rect 7060 4863 7376 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 2479 4384 2795 4385
rect 2479 4320 2485 4384
rect 2549 4320 2565 4384
rect 2629 4320 2645 4384
rect 2709 4320 2725 4384
rect 2789 4320 2795 4384
rect 2479 4319 2795 4320
rect 4226 4384 4542 4385
rect 4226 4320 4232 4384
rect 4296 4320 4312 4384
rect 4376 4320 4392 4384
rect 4456 4320 4472 4384
rect 4536 4320 4542 4384
rect 4226 4319 4542 4320
rect 5973 4384 6289 4385
rect 5973 4320 5979 4384
rect 6043 4320 6059 4384
rect 6123 4320 6139 4384
rect 6203 4320 6219 4384
rect 6283 4320 6289 4384
rect 5973 4319 6289 4320
rect 7720 4384 8036 4385
rect 7720 4320 7726 4384
rect 7790 4320 7806 4384
rect 7870 4320 7886 4384
rect 7950 4320 7966 4384
rect 8030 4320 8036 4384
rect 7720 4319 8036 4320
rect 8109 4178 8175 4181
rect 8404 4178 9204 4208
rect 8109 4176 9204 4178
rect 8109 4120 8114 4176
rect 8170 4120 9204 4176
rect 8109 4118 9204 4120
rect 8109 4115 8175 4118
rect 8404 4088 9204 4118
rect 3509 4042 3575 4045
rect 2730 4040 3575 4042
rect 2730 3984 3514 4040
rect 3570 3984 3575 4040
rect 2730 3982 3575 3984
rect 1819 3840 2135 3841
rect 1819 3776 1825 3840
rect 1889 3776 1905 3840
rect 1969 3776 1985 3840
rect 2049 3776 2065 3840
rect 2129 3776 2135 3840
rect 1819 3775 2135 3776
rect 0 3498 800 3528
rect 2730 3498 2790 3982
rect 3509 3979 3575 3982
rect 3566 3840 3882 3841
rect 3566 3776 3572 3840
rect 3636 3776 3652 3840
rect 3716 3776 3732 3840
rect 3796 3776 3812 3840
rect 3876 3776 3882 3840
rect 3566 3775 3882 3776
rect 5313 3840 5629 3841
rect 5313 3776 5319 3840
rect 5383 3776 5399 3840
rect 5463 3776 5479 3840
rect 5543 3776 5559 3840
rect 5623 3776 5629 3840
rect 5313 3775 5629 3776
rect 7060 3840 7376 3841
rect 7060 3776 7066 3840
rect 7130 3776 7146 3840
rect 7210 3776 7226 3840
rect 7290 3776 7306 3840
rect 7370 3776 7376 3840
rect 7060 3775 7376 3776
rect 0 3438 2790 3498
rect 0 3408 800 3438
rect 2479 3296 2795 3297
rect 2479 3232 2485 3296
rect 2549 3232 2565 3296
rect 2629 3232 2645 3296
rect 2709 3232 2725 3296
rect 2789 3232 2795 3296
rect 2479 3231 2795 3232
rect 4226 3296 4542 3297
rect 4226 3232 4232 3296
rect 4296 3232 4312 3296
rect 4376 3232 4392 3296
rect 4456 3232 4472 3296
rect 4536 3232 4542 3296
rect 4226 3231 4542 3232
rect 5973 3296 6289 3297
rect 5973 3232 5979 3296
rect 6043 3232 6059 3296
rect 6123 3232 6139 3296
rect 6203 3232 6219 3296
rect 6283 3232 6289 3296
rect 5973 3231 6289 3232
rect 7720 3296 8036 3297
rect 7720 3232 7726 3296
rect 7790 3232 7806 3296
rect 7870 3232 7886 3296
rect 7950 3232 7966 3296
rect 8030 3232 8036 3296
rect 7720 3231 8036 3232
rect 2129 2954 2195 2957
rect 2998 2954 3004 2956
rect 2129 2952 3004 2954
rect 2129 2896 2134 2952
rect 2190 2896 3004 2952
rect 2129 2894 3004 2896
rect 2129 2891 2195 2894
rect 2998 2892 3004 2894
rect 3068 2954 3074 2956
rect 5809 2954 5875 2957
rect 3068 2952 5875 2954
rect 3068 2896 5814 2952
rect 5870 2896 5875 2952
rect 3068 2894 5875 2896
rect 3068 2892 3074 2894
rect 5809 2891 5875 2894
rect 1819 2752 2135 2753
rect 1819 2688 1825 2752
rect 1889 2688 1905 2752
rect 1969 2688 1985 2752
rect 2049 2688 2065 2752
rect 2129 2688 2135 2752
rect 1819 2687 2135 2688
rect 3566 2752 3882 2753
rect 3566 2688 3572 2752
rect 3636 2688 3652 2752
rect 3716 2688 3732 2752
rect 3796 2688 3812 2752
rect 3876 2688 3882 2752
rect 3566 2687 3882 2688
rect 5313 2752 5629 2753
rect 5313 2688 5319 2752
rect 5383 2688 5399 2752
rect 5463 2688 5479 2752
rect 5543 2688 5559 2752
rect 5623 2688 5629 2752
rect 5313 2687 5629 2688
rect 7060 2752 7376 2753
rect 7060 2688 7066 2752
rect 7130 2688 7146 2752
rect 7210 2688 7226 2752
rect 7290 2688 7306 2752
rect 7370 2688 7376 2752
rect 7060 2687 7376 2688
rect 4889 2410 4955 2413
rect 4889 2408 8218 2410
rect 4889 2352 4894 2408
rect 4950 2352 8218 2408
rect 4889 2350 8218 2352
rect 4889 2347 4955 2350
rect 2479 2208 2795 2209
rect 2479 2144 2485 2208
rect 2549 2144 2565 2208
rect 2629 2144 2645 2208
rect 2709 2144 2725 2208
rect 2789 2144 2795 2208
rect 2479 2143 2795 2144
rect 4226 2208 4542 2209
rect 4226 2144 4232 2208
rect 4296 2144 4312 2208
rect 4376 2144 4392 2208
rect 4456 2144 4472 2208
rect 4536 2144 4542 2208
rect 4226 2143 4542 2144
rect 5973 2208 6289 2209
rect 5973 2144 5979 2208
rect 6043 2144 6059 2208
rect 6123 2144 6139 2208
rect 6203 2144 6219 2208
rect 6283 2144 6289 2208
rect 5973 2143 6289 2144
rect 7720 2208 8036 2209
rect 7720 2144 7726 2208
rect 7790 2144 7806 2208
rect 7870 2144 7886 2208
rect 7950 2144 7966 2208
rect 8030 2144 8036 2208
rect 7720 2143 8036 2144
rect 8158 2138 8218 2350
rect 8404 2138 9204 2168
rect 8158 2078 9204 2138
rect 8404 2048 9204 2078
rect 0 1458 800 1488
rect 3141 1458 3207 1461
rect 0 1456 3207 1458
rect 0 1400 3146 1456
rect 3202 1400 3207 1456
rect 0 1398 3207 1400
rect 0 1368 800 1398
rect 3141 1395 3207 1398
rect 2262 716 2268 780
rect 2332 778 2338 780
rect 3325 778 3391 781
rect 2332 776 3391 778
rect 2332 720 3330 776
rect 3386 720 3391 776
rect 2332 718 3391 720
rect 2332 716 2338 718
rect 3325 715 3391 718
rect 4153 778 4219 781
rect 8404 778 9204 808
rect 4153 776 9204 778
rect 4153 720 4158 776
rect 4214 720 9204 776
rect 4153 718 9204 720
rect 4153 715 4219 718
rect 8404 688 9204 718
<< via3 >>
rect 2485 8732 2549 8736
rect 2485 8676 2489 8732
rect 2489 8676 2545 8732
rect 2545 8676 2549 8732
rect 2485 8672 2549 8676
rect 2565 8732 2629 8736
rect 2565 8676 2569 8732
rect 2569 8676 2625 8732
rect 2625 8676 2629 8732
rect 2565 8672 2629 8676
rect 2645 8732 2709 8736
rect 2645 8676 2649 8732
rect 2649 8676 2705 8732
rect 2705 8676 2709 8732
rect 2645 8672 2709 8676
rect 2725 8732 2789 8736
rect 2725 8676 2729 8732
rect 2729 8676 2785 8732
rect 2785 8676 2789 8732
rect 2725 8672 2789 8676
rect 4232 8732 4296 8736
rect 4232 8676 4236 8732
rect 4236 8676 4292 8732
rect 4292 8676 4296 8732
rect 4232 8672 4296 8676
rect 4312 8732 4376 8736
rect 4312 8676 4316 8732
rect 4316 8676 4372 8732
rect 4372 8676 4376 8732
rect 4312 8672 4376 8676
rect 4392 8732 4456 8736
rect 4392 8676 4396 8732
rect 4396 8676 4452 8732
rect 4452 8676 4456 8732
rect 4392 8672 4456 8676
rect 4472 8732 4536 8736
rect 4472 8676 4476 8732
rect 4476 8676 4532 8732
rect 4532 8676 4536 8732
rect 4472 8672 4536 8676
rect 5979 8732 6043 8736
rect 5979 8676 5983 8732
rect 5983 8676 6039 8732
rect 6039 8676 6043 8732
rect 5979 8672 6043 8676
rect 6059 8732 6123 8736
rect 6059 8676 6063 8732
rect 6063 8676 6119 8732
rect 6119 8676 6123 8732
rect 6059 8672 6123 8676
rect 6139 8732 6203 8736
rect 6139 8676 6143 8732
rect 6143 8676 6199 8732
rect 6199 8676 6203 8732
rect 6139 8672 6203 8676
rect 6219 8732 6283 8736
rect 6219 8676 6223 8732
rect 6223 8676 6279 8732
rect 6279 8676 6283 8732
rect 6219 8672 6283 8676
rect 7726 8732 7790 8736
rect 7726 8676 7730 8732
rect 7730 8676 7786 8732
rect 7786 8676 7790 8732
rect 7726 8672 7790 8676
rect 7806 8732 7870 8736
rect 7806 8676 7810 8732
rect 7810 8676 7866 8732
rect 7866 8676 7870 8732
rect 7806 8672 7870 8676
rect 7886 8732 7950 8736
rect 7886 8676 7890 8732
rect 7890 8676 7946 8732
rect 7946 8676 7950 8732
rect 7886 8672 7950 8676
rect 7966 8732 8030 8736
rect 7966 8676 7970 8732
rect 7970 8676 8026 8732
rect 8026 8676 8030 8732
rect 7966 8672 8030 8676
rect 1825 8188 1889 8192
rect 1825 8132 1829 8188
rect 1829 8132 1885 8188
rect 1885 8132 1889 8188
rect 1825 8128 1889 8132
rect 1905 8188 1969 8192
rect 1905 8132 1909 8188
rect 1909 8132 1965 8188
rect 1965 8132 1969 8188
rect 1905 8128 1969 8132
rect 1985 8188 2049 8192
rect 1985 8132 1989 8188
rect 1989 8132 2045 8188
rect 2045 8132 2049 8188
rect 1985 8128 2049 8132
rect 2065 8188 2129 8192
rect 2065 8132 2069 8188
rect 2069 8132 2125 8188
rect 2125 8132 2129 8188
rect 2065 8128 2129 8132
rect 3572 8188 3636 8192
rect 3572 8132 3576 8188
rect 3576 8132 3632 8188
rect 3632 8132 3636 8188
rect 3572 8128 3636 8132
rect 3652 8188 3716 8192
rect 3652 8132 3656 8188
rect 3656 8132 3712 8188
rect 3712 8132 3716 8188
rect 3652 8128 3716 8132
rect 3732 8188 3796 8192
rect 3732 8132 3736 8188
rect 3736 8132 3792 8188
rect 3792 8132 3796 8188
rect 3732 8128 3796 8132
rect 3812 8188 3876 8192
rect 3812 8132 3816 8188
rect 3816 8132 3872 8188
rect 3872 8132 3876 8188
rect 3812 8128 3876 8132
rect 5319 8188 5383 8192
rect 5319 8132 5323 8188
rect 5323 8132 5379 8188
rect 5379 8132 5383 8188
rect 5319 8128 5383 8132
rect 5399 8188 5463 8192
rect 5399 8132 5403 8188
rect 5403 8132 5459 8188
rect 5459 8132 5463 8188
rect 5399 8128 5463 8132
rect 5479 8188 5543 8192
rect 5479 8132 5483 8188
rect 5483 8132 5539 8188
rect 5539 8132 5543 8188
rect 5479 8128 5543 8132
rect 5559 8188 5623 8192
rect 5559 8132 5563 8188
rect 5563 8132 5619 8188
rect 5619 8132 5623 8188
rect 5559 8128 5623 8132
rect 7066 8188 7130 8192
rect 7066 8132 7070 8188
rect 7070 8132 7126 8188
rect 7126 8132 7130 8188
rect 7066 8128 7130 8132
rect 7146 8188 7210 8192
rect 7146 8132 7150 8188
rect 7150 8132 7206 8188
rect 7206 8132 7210 8188
rect 7146 8128 7210 8132
rect 7226 8188 7290 8192
rect 7226 8132 7230 8188
rect 7230 8132 7286 8188
rect 7286 8132 7290 8188
rect 7226 8128 7290 8132
rect 7306 8188 7370 8192
rect 7306 8132 7310 8188
rect 7310 8132 7366 8188
rect 7366 8132 7370 8188
rect 7306 8128 7370 8132
rect 2485 7644 2549 7648
rect 2485 7588 2489 7644
rect 2489 7588 2545 7644
rect 2545 7588 2549 7644
rect 2485 7584 2549 7588
rect 2565 7644 2629 7648
rect 2565 7588 2569 7644
rect 2569 7588 2625 7644
rect 2625 7588 2629 7644
rect 2565 7584 2629 7588
rect 2645 7644 2709 7648
rect 2645 7588 2649 7644
rect 2649 7588 2705 7644
rect 2705 7588 2709 7644
rect 2645 7584 2709 7588
rect 2725 7644 2789 7648
rect 2725 7588 2729 7644
rect 2729 7588 2785 7644
rect 2785 7588 2789 7644
rect 2725 7584 2789 7588
rect 4232 7644 4296 7648
rect 4232 7588 4236 7644
rect 4236 7588 4292 7644
rect 4292 7588 4296 7644
rect 4232 7584 4296 7588
rect 4312 7644 4376 7648
rect 4312 7588 4316 7644
rect 4316 7588 4372 7644
rect 4372 7588 4376 7644
rect 4312 7584 4376 7588
rect 4392 7644 4456 7648
rect 4392 7588 4396 7644
rect 4396 7588 4452 7644
rect 4452 7588 4456 7644
rect 4392 7584 4456 7588
rect 4472 7644 4536 7648
rect 4472 7588 4476 7644
rect 4476 7588 4532 7644
rect 4532 7588 4536 7644
rect 4472 7584 4536 7588
rect 5979 7644 6043 7648
rect 5979 7588 5983 7644
rect 5983 7588 6039 7644
rect 6039 7588 6043 7644
rect 5979 7584 6043 7588
rect 6059 7644 6123 7648
rect 6059 7588 6063 7644
rect 6063 7588 6119 7644
rect 6119 7588 6123 7644
rect 6059 7584 6123 7588
rect 6139 7644 6203 7648
rect 6139 7588 6143 7644
rect 6143 7588 6199 7644
rect 6199 7588 6203 7644
rect 6139 7584 6203 7588
rect 6219 7644 6283 7648
rect 6219 7588 6223 7644
rect 6223 7588 6279 7644
rect 6279 7588 6283 7644
rect 6219 7584 6283 7588
rect 7726 7644 7790 7648
rect 7726 7588 7730 7644
rect 7730 7588 7786 7644
rect 7786 7588 7790 7644
rect 7726 7584 7790 7588
rect 7806 7644 7870 7648
rect 7806 7588 7810 7644
rect 7810 7588 7866 7644
rect 7866 7588 7870 7644
rect 7806 7584 7870 7588
rect 7886 7644 7950 7648
rect 7886 7588 7890 7644
rect 7890 7588 7946 7644
rect 7946 7588 7950 7644
rect 7886 7584 7950 7588
rect 7966 7644 8030 7648
rect 7966 7588 7970 7644
rect 7970 7588 8026 7644
rect 8026 7588 8030 7644
rect 7966 7584 8030 7588
rect 1825 7100 1889 7104
rect 1825 7044 1829 7100
rect 1829 7044 1885 7100
rect 1885 7044 1889 7100
rect 1825 7040 1889 7044
rect 1905 7100 1969 7104
rect 1905 7044 1909 7100
rect 1909 7044 1965 7100
rect 1965 7044 1969 7100
rect 1905 7040 1969 7044
rect 1985 7100 2049 7104
rect 1985 7044 1989 7100
rect 1989 7044 2045 7100
rect 2045 7044 2049 7100
rect 1985 7040 2049 7044
rect 2065 7100 2129 7104
rect 2065 7044 2069 7100
rect 2069 7044 2125 7100
rect 2125 7044 2129 7100
rect 2065 7040 2129 7044
rect 3572 7100 3636 7104
rect 3572 7044 3576 7100
rect 3576 7044 3632 7100
rect 3632 7044 3636 7100
rect 3572 7040 3636 7044
rect 3652 7100 3716 7104
rect 3652 7044 3656 7100
rect 3656 7044 3712 7100
rect 3712 7044 3716 7100
rect 3652 7040 3716 7044
rect 3732 7100 3796 7104
rect 3732 7044 3736 7100
rect 3736 7044 3792 7100
rect 3792 7044 3796 7100
rect 3732 7040 3796 7044
rect 3812 7100 3876 7104
rect 3812 7044 3816 7100
rect 3816 7044 3872 7100
rect 3872 7044 3876 7100
rect 3812 7040 3876 7044
rect 5319 7100 5383 7104
rect 5319 7044 5323 7100
rect 5323 7044 5379 7100
rect 5379 7044 5383 7100
rect 5319 7040 5383 7044
rect 5399 7100 5463 7104
rect 5399 7044 5403 7100
rect 5403 7044 5459 7100
rect 5459 7044 5463 7100
rect 5399 7040 5463 7044
rect 5479 7100 5543 7104
rect 5479 7044 5483 7100
rect 5483 7044 5539 7100
rect 5539 7044 5543 7100
rect 5479 7040 5543 7044
rect 5559 7100 5623 7104
rect 5559 7044 5563 7100
rect 5563 7044 5619 7100
rect 5619 7044 5623 7100
rect 5559 7040 5623 7044
rect 7066 7100 7130 7104
rect 7066 7044 7070 7100
rect 7070 7044 7126 7100
rect 7126 7044 7130 7100
rect 7066 7040 7130 7044
rect 7146 7100 7210 7104
rect 7146 7044 7150 7100
rect 7150 7044 7206 7100
rect 7206 7044 7210 7100
rect 7146 7040 7210 7044
rect 7226 7100 7290 7104
rect 7226 7044 7230 7100
rect 7230 7044 7286 7100
rect 7286 7044 7290 7100
rect 7226 7040 7290 7044
rect 7306 7100 7370 7104
rect 7306 7044 7310 7100
rect 7310 7044 7366 7100
rect 7366 7044 7370 7100
rect 7306 7040 7370 7044
rect 2485 6556 2549 6560
rect 2485 6500 2489 6556
rect 2489 6500 2545 6556
rect 2545 6500 2549 6556
rect 2485 6496 2549 6500
rect 2565 6556 2629 6560
rect 2565 6500 2569 6556
rect 2569 6500 2625 6556
rect 2625 6500 2629 6556
rect 2565 6496 2629 6500
rect 2645 6556 2709 6560
rect 2645 6500 2649 6556
rect 2649 6500 2705 6556
rect 2705 6500 2709 6556
rect 2645 6496 2709 6500
rect 2725 6556 2789 6560
rect 2725 6500 2729 6556
rect 2729 6500 2785 6556
rect 2785 6500 2789 6556
rect 2725 6496 2789 6500
rect 4232 6556 4296 6560
rect 4232 6500 4236 6556
rect 4236 6500 4292 6556
rect 4292 6500 4296 6556
rect 4232 6496 4296 6500
rect 4312 6556 4376 6560
rect 4312 6500 4316 6556
rect 4316 6500 4372 6556
rect 4372 6500 4376 6556
rect 4312 6496 4376 6500
rect 4392 6556 4456 6560
rect 4392 6500 4396 6556
rect 4396 6500 4452 6556
rect 4452 6500 4456 6556
rect 4392 6496 4456 6500
rect 4472 6556 4536 6560
rect 4472 6500 4476 6556
rect 4476 6500 4532 6556
rect 4532 6500 4536 6556
rect 4472 6496 4536 6500
rect 5979 6556 6043 6560
rect 5979 6500 5983 6556
rect 5983 6500 6039 6556
rect 6039 6500 6043 6556
rect 5979 6496 6043 6500
rect 6059 6556 6123 6560
rect 6059 6500 6063 6556
rect 6063 6500 6119 6556
rect 6119 6500 6123 6556
rect 6059 6496 6123 6500
rect 6139 6556 6203 6560
rect 6139 6500 6143 6556
rect 6143 6500 6199 6556
rect 6199 6500 6203 6556
rect 6139 6496 6203 6500
rect 6219 6556 6283 6560
rect 6219 6500 6223 6556
rect 6223 6500 6279 6556
rect 6279 6500 6283 6556
rect 6219 6496 6283 6500
rect 7726 6556 7790 6560
rect 7726 6500 7730 6556
rect 7730 6500 7786 6556
rect 7786 6500 7790 6556
rect 7726 6496 7790 6500
rect 7806 6556 7870 6560
rect 7806 6500 7810 6556
rect 7810 6500 7866 6556
rect 7866 6500 7870 6556
rect 7806 6496 7870 6500
rect 7886 6556 7950 6560
rect 7886 6500 7890 6556
rect 7890 6500 7946 6556
rect 7946 6500 7950 6556
rect 7886 6496 7950 6500
rect 7966 6556 8030 6560
rect 7966 6500 7970 6556
rect 7970 6500 8026 6556
rect 8026 6500 8030 6556
rect 7966 6496 8030 6500
rect 2268 6352 2332 6356
rect 2268 6296 2282 6352
rect 2282 6296 2332 6352
rect 2268 6292 2332 6296
rect 1825 6012 1889 6016
rect 1825 5956 1829 6012
rect 1829 5956 1885 6012
rect 1885 5956 1889 6012
rect 1825 5952 1889 5956
rect 1905 6012 1969 6016
rect 1905 5956 1909 6012
rect 1909 5956 1965 6012
rect 1965 5956 1969 6012
rect 1905 5952 1969 5956
rect 1985 6012 2049 6016
rect 1985 5956 1989 6012
rect 1989 5956 2045 6012
rect 2045 5956 2049 6012
rect 1985 5952 2049 5956
rect 2065 6012 2129 6016
rect 2065 5956 2069 6012
rect 2069 5956 2125 6012
rect 2125 5956 2129 6012
rect 2065 5952 2129 5956
rect 3572 6012 3636 6016
rect 3572 5956 3576 6012
rect 3576 5956 3632 6012
rect 3632 5956 3636 6012
rect 3572 5952 3636 5956
rect 3652 6012 3716 6016
rect 3652 5956 3656 6012
rect 3656 5956 3712 6012
rect 3712 5956 3716 6012
rect 3652 5952 3716 5956
rect 3732 6012 3796 6016
rect 3732 5956 3736 6012
rect 3736 5956 3792 6012
rect 3792 5956 3796 6012
rect 3732 5952 3796 5956
rect 3812 6012 3876 6016
rect 3812 5956 3816 6012
rect 3816 5956 3872 6012
rect 3872 5956 3876 6012
rect 3812 5952 3876 5956
rect 5319 6012 5383 6016
rect 5319 5956 5323 6012
rect 5323 5956 5379 6012
rect 5379 5956 5383 6012
rect 5319 5952 5383 5956
rect 5399 6012 5463 6016
rect 5399 5956 5403 6012
rect 5403 5956 5459 6012
rect 5459 5956 5463 6012
rect 5399 5952 5463 5956
rect 5479 6012 5543 6016
rect 5479 5956 5483 6012
rect 5483 5956 5539 6012
rect 5539 5956 5543 6012
rect 5479 5952 5543 5956
rect 5559 6012 5623 6016
rect 5559 5956 5563 6012
rect 5563 5956 5619 6012
rect 5619 5956 5623 6012
rect 5559 5952 5623 5956
rect 7066 6012 7130 6016
rect 7066 5956 7070 6012
rect 7070 5956 7126 6012
rect 7126 5956 7130 6012
rect 7066 5952 7130 5956
rect 7146 6012 7210 6016
rect 7146 5956 7150 6012
rect 7150 5956 7206 6012
rect 7206 5956 7210 6012
rect 7146 5952 7210 5956
rect 7226 6012 7290 6016
rect 7226 5956 7230 6012
rect 7230 5956 7286 6012
rect 7286 5956 7290 6012
rect 7226 5952 7290 5956
rect 7306 6012 7370 6016
rect 7306 5956 7310 6012
rect 7310 5956 7366 6012
rect 7366 5956 7370 6012
rect 7306 5952 7370 5956
rect 2485 5468 2549 5472
rect 2485 5412 2489 5468
rect 2489 5412 2545 5468
rect 2545 5412 2549 5468
rect 2485 5408 2549 5412
rect 2565 5468 2629 5472
rect 2565 5412 2569 5468
rect 2569 5412 2625 5468
rect 2625 5412 2629 5468
rect 2565 5408 2629 5412
rect 2645 5468 2709 5472
rect 2645 5412 2649 5468
rect 2649 5412 2705 5468
rect 2705 5412 2709 5468
rect 2645 5408 2709 5412
rect 2725 5468 2789 5472
rect 2725 5412 2729 5468
rect 2729 5412 2785 5468
rect 2785 5412 2789 5468
rect 2725 5408 2789 5412
rect 4232 5468 4296 5472
rect 4232 5412 4236 5468
rect 4236 5412 4292 5468
rect 4292 5412 4296 5468
rect 4232 5408 4296 5412
rect 4312 5468 4376 5472
rect 4312 5412 4316 5468
rect 4316 5412 4372 5468
rect 4372 5412 4376 5468
rect 4312 5408 4376 5412
rect 4392 5468 4456 5472
rect 4392 5412 4396 5468
rect 4396 5412 4452 5468
rect 4452 5412 4456 5468
rect 4392 5408 4456 5412
rect 4472 5468 4536 5472
rect 4472 5412 4476 5468
rect 4476 5412 4532 5468
rect 4532 5412 4536 5468
rect 4472 5408 4536 5412
rect 5979 5468 6043 5472
rect 5979 5412 5983 5468
rect 5983 5412 6039 5468
rect 6039 5412 6043 5468
rect 5979 5408 6043 5412
rect 6059 5468 6123 5472
rect 6059 5412 6063 5468
rect 6063 5412 6119 5468
rect 6119 5412 6123 5468
rect 6059 5408 6123 5412
rect 6139 5468 6203 5472
rect 6139 5412 6143 5468
rect 6143 5412 6199 5468
rect 6199 5412 6203 5468
rect 6139 5408 6203 5412
rect 6219 5468 6283 5472
rect 6219 5412 6223 5468
rect 6223 5412 6279 5468
rect 6279 5412 6283 5468
rect 6219 5408 6283 5412
rect 7726 5468 7790 5472
rect 7726 5412 7730 5468
rect 7730 5412 7786 5468
rect 7786 5412 7790 5468
rect 7726 5408 7790 5412
rect 7806 5468 7870 5472
rect 7806 5412 7810 5468
rect 7810 5412 7866 5468
rect 7866 5412 7870 5468
rect 7806 5408 7870 5412
rect 7886 5468 7950 5472
rect 7886 5412 7890 5468
rect 7890 5412 7946 5468
rect 7946 5412 7950 5468
rect 7886 5408 7950 5412
rect 7966 5468 8030 5472
rect 7966 5412 7970 5468
rect 7970 5412 8026 5468
rect 8026 5412 8030 5468
rect 7966 5408 8030 5412
rect 3004 5068 3068 5132
rect 1825 4924 1889 4928
rect 1825 4868 1829 4924
rect 1829 4868 1885 4924
rect 1885 4868 1889 4924
rect 1825 4864 1889 4868
rect 1905 4924 1969 4928
rect 1905 4868 1909 4924
rect 1909 4868 1965 4924
rect 1965 4868 1969 4924
rect 1905 4864 1969 4868
rect 1985 4924 2049 4928
rect 1985 4868 1989 4924
rect 1989 4868 2045 4924
rect 2045 4868 2049 4924
rect 1985 4864 2049 4868
rect 2065 4924 2129 4928
rect 2065 4868 2069 4924
rect 2069 4868 2125 4924
rect 2125 4868 2129 4924
rect 2065 4864 2129 4868
rect 3572 4924 3636 4928
rect 3572 4868 3576 4924
rect 3576 4868 3632 4924
rect 3632 4868 3636 4924
rect 3572 4864 3636 4868
rect 3652 4924 3716 4928
rect 3652 4868 3656 4924
rect 3656 4868 3712 4924
rect 3712 4868 3716 4924
rect 3652 4864 3716 4868
rect 3732 4924 3796 4928
rect 3732 4868 3736 4924
rect 3736 4868 3792 4924
rect 3792 4868 3796 4924
rect 3732 4864 3796 4868
rect 3812 4924 3876 4928
rect 3812 4868 3816 4924
rect 3816 4868 3872 4924
rect 3872 4868 3876 4924
rect 3812 4864 3876 4868
rect 5319 4924 5383 4928
rect 5319 4868 5323 4924
rect 5323 4868 5379 4924
rect 5379 4868 5383 4924
rect 5319 4864 5383 4868
rect 5399 4924 5463 4928
rect 5399 4868 5403 4924
rect 5403 4868 5459 4924
rect 5459 4868 5463 4924
rect 5399 4864 5463 4868
rect 5479 4924 5543 4928
rect 5479 4868 5483 4924
rect 5483 4868 5539 4924
rect 5539 4868 5543 4924
rect 5479 4864 5543 4868
rect 5559 4924 5623 4928
rect 5559 4868 5563 4924
rect 5563 4868 5619 4924
rect 5619 4868 5623 4924
rect 5559 4864 5623 4868
rect 7066 4924 7130 4928
rect 7066 4868 7070 4924
rect 7070 4868 7126 4924
rect 7126 4868 7130 4924
rect 7066 4864 7130 4868
rect 7146 4924 7210 4928
rect 7146 4868 7150 4924
rect 7150 4868 7206 4924
rect 7206 4868 7210 4924
rect 7146 4864 7210 4868
rect 7226 4924 7290 4928
rect 7226 4868 7230 4924
rect 7230 4868 7286 4924
rect 7286 4868 7290 4924
rect 7226 4864 7290 4868
rect 7306 4924 7370 4928
rect 7306 4868 7310 4924
rect 7310 4868 7366 4924
rect 7366 4868 7370 4924
rect 7306 4864 7370 4868
rect 2485 4380 2549 4384
rect 2485 4324 2489 4380
rect 2489 4324 2545 4380
rect 2545 4324 2549 4380
rect 2485 4320 2549 4324
rect 2565 4380 2629 4384
rect 2565 4324 2569 4380
rect 2569 4324 2625 4380
rect 2625 4324 2629 4380
rect 2565 4320 2629 4324
rect 2645 4380 2709 4384
rect 2645 4324 2649 4380
rect 2649 4324 2705 4380
rect 2705 4324 2709 4380
rect 2645 4320 2709 4324
rect 2725 4380 2789 4384
rect 2725 4324 2729 4380
rect 2729 4324 2785 4380
rect 2785 4324 2789 4380
rect 2725 4320 2789 4324
rect 4232 4380 4296 4384
rect 4232 4324 4236 4380
rect 4236 4324 4292 4380
rect 4292 4324 4296 4380
rect 4232 4320 4296 4324
rect 4312 4380 4376 4384
rect 4312 4324 4316 4380
rect 4316 4324 4372 4380
rect 4372 4324 4376 4380
rect 4312 4320 4376 4324
rect 4392 4380 4456 4384
rect 4392 4324 4396 4380
rect 4396 4324 4452 4380
rect 4452 4324 4456 4380
rect 4392 4320 4456 4324
rect 4472 4380 4536 4384
rect 4472 4324 4476 4380
rect 4476 4324 4532 4380
rect 4532 4324 4536 4380
rect 4472 4320 4536 4324
rect 5979 4380 6043 4384
rect 5979 4324 5983 4380
rect 5983 4324 6039 4380
rect 6039 4324 6043 4380
rect 5979 4320 6043 4324
rect 6059 4380 6123 4384
rect 6059 4324 6063 4380
rect 6063 4324 6119 4380
rect 6119 4324 6123 4380
rect 6059 4320 6123 4324
rect 6139 4380 6203 4384
rect 6139 4324 6143 4380
rect 6143 4324 6199 4380
rect 6199 4324 6203 4380
rect 6139 4320 6203 4324
rect 6219 4380 6283 4384
rect 6219 4324 6223 4380
rect 6223 4324 6279 4380
rect 6279 4324 6283 4380
rect 6219 4320 6283 4324
rect 7726 4380 7790 4384
rect 7726 4324 7730 4380
rect 7730 4324 7786 4380
rect 7786 4324 7790 4380
rect 7726 4320 7790 4324
rect 7806 4380 7870 4384
rect 7806 4324 7810 4380
rect 7810 4324 7866 4380
rect 7866 4324 7870 4380
rect 7806 4320 7870 4324
rect 7886 4380 7950 4384
rect 7886 4324 7890 4380
rect 7890 4324 7946 4380
rect 7946 4324 7950 4380
rect 7886 4320 7950 4324
rect 7966 4380 8030 4384
rect 7966 4324 7970 4380
rect 7970 4324 8026 4380
rect 8026 4324 8030 4380
rect 7966 4320 8030 4324
rect 1825 3836 1889 3840
rect 1825 3780 1829 3836
rect 1829 3780 1885 3836
rect 1885 3780 1889 3836
rect 1825 3776 1889 3780
rect 1905 3836 1969 3840
rect 1905 3780 1909 3836
rect 1909 3780 1965 3836
rect 1965 3780 1969 3836
rect 1905 3776 1969 3780
rect 1985 3836 2049 3840
rect 1985 3780 1989 3836
rect 1989 3780 2045 3836
rect 2045 3780 2049 3836
rect 1985 3776 2049 3780
rect 2065 3836 2129 3840
rect 2065 3780 2069 3836
rect 2069 3780 2125 3836
rect 2125 3780 2129 3836
rect 2065 3776 2129 3780
rect 3572 3836 3636 3840
rect 3572 3780 3576 3836
rect 3576 3780 3632 3836
rect 3632 3780 3636 3836
rect 3572 3776 3636 3780
rect 3652 3836 3716 3840
rect 3652 3780 3656 3836
rect 3656 3780 3712 3836
rect 3712 3780 3716 3836
rect 3652 3776 3716 3780
rect 3732 3836 3796 3840
rect 3732 3780 3736 3836
rect 3736 3780 3792 3836
rect 3792 3780 3796 3836
rect 3732 3776 3796 3780
rect 3812 3836 3876 3840
rect 3812 3780 3816 3836
rect 3816 3780 3872 3836
rect 3872 3780 3876 3836
rect 3812 3776 3876 3780
rect 5319 3836 5383 3840
rect 5319 3780 5323 3836
rect 5323 3780 5379 3836
rect 5379 3780 5383 3836
rect 5319 3776 5383 3780
rect 5399 3836 5463 3840
rect 5399 3780 5403 3836
rect 5403 3780 5459 3836
rect 5459 3780 5463 3836
rect 5399 3776 5463 3780
rect 5479 3836 5543 3840
rect 5479 3780 5483 3836
rect 5483 3780 5539 3836
rect 5539 3780 5543 3836
rect 5479 3776 5543 3780
rect 5559 3836 5623 3840
rect 5559 3780 5563 3836
rect 5563 3780 5619 3836
rect 5619 3780 5623 3836
rect 5559 3776 5623 3780
rect 7066 3836 7130 3840
rect 7066 3780 7070 3836
rect 7070 3780 7126 3836
rect 7126 3780 7130 3836
rect 7066 3776 7130 3780
rect 7146 3836 7210 3840
rect 7146 3780 7150 3836
rect 7150 3780 7206 3836
rect 7206 3780 7210 3836
rect 7146 3776 7210 3780
rect 7226 3836 7290 3840
rect 7226 3780 7230 3836
rect 7230 3780 7286 3836
rect 7286 3780 7290 3836
rect 7226 3776 7290 3780
rect 7306 3836 7370 3840
rect 7306 3780 7310 3836
rect 7310 3780 7366 3836
rect 7366 3780 7370 3836
rect 7306 3776 7370 3780
rect 2485 3292 2549 3296
rect 2485 3236 2489 3292
rect 2489 3236 2545 3292
rect 2545 3236 2549 3292
rect 2485 3232 2549 3236
rect 2565 3292 2629 3296
rect 2565 3236 2569 3292
rect 2569 3236 2625 3292
rect 2625 3236 2629 3292
rect 2565 3232 2629 3236
rect 2645 3292 2709 3296
rect 2645 3236 2649 3292
rect 2649 3236 2705 3292
rect 2705 3236 2709 3292
rect 2645 3232 2709 3236
rect 2725 3292 2789 3296
rect 2725 3236 2729 3292
rect 2729 3236 2785 3292
rect 2785 3236 2789 3292
rect 2725 3232 2789 3236
rect 4232 3292 4296 3296
rect 4232 3236 4236 3292
rect 4236 3236 4292 3292
rect 4292 3236 4296 3292
rect 4232 3232 4296 3236
rect 4312 3292 4376 3296
rect 4312 3236 4316 3292
rect 4316 3236 4372 3292
rect 4372 3236 4376 3292
rect 4312 3232 4376 3236
rect 4392 3292 4456 3296
rect 4392 3236 4396 3292
rect 4396 3236 4452 3292
rect 4452 3236 4456 3292
rect 4392 3232 4456 3236
rect 4472 3292 4536 3296
rect 4472 3236 4476 3292
rect 4476 3236 4532 3292
rect 4532 3236 4536 3292
rect 4472 3232 4536 3236
rect 5979 3292 6043 3296
rect 5979 3236 5983 3292
rect 5983 3236 6039 3292
rect 6039 3236 6043 3292
rect 5979 3232 6043 3236
rect 6059 3292 6123 3296
rect 6059 3236 6063 3292
rect 6063 3236 6119 3292
rect 6119 3236 6123 3292
rect 6059 3232 6123 3236
rect 6139 3292 6203 3296
rect 6139 3236 6143 3292
rect 6143 3236 6199 3292
rect 6199 3236 6203 3292
rect 6139 3232 6203 3236
rect 6219 3292 6283 3296
rect 6219 3236 6223 3292
rect 6223 3236 6279 3292
rect 6279 3236 6283 3292
rect 6219 3232 6283 3236
rect 7726 3292 7790 3296
rect 7726 3236 7730 3292
rect 7730 3236 7786 3292
rect 7786 3236 7790 3292
rect 7726 3232 7790 3236
rect 7806 3292 7870 3296
rect 7806 3236 7810 3292
rect 7810 3236 7866 3292
rect 7866 3236 7870 3292
rect 7806 3232 7870 3236
rect 7886 3292 7950 3296
rect 7886 3236 7890 3292
rect 7890 3236 7946 3292
rect 7946 3236 7950 3292
rect 7886 3232 7950 3236
rect 7966 3292 8030 3296
rect 7966 3236 7970 3292
rect 7970 3236 8026 3292
rect 8026 3236 8030 3292
rect 7966 3232 8030 3236
rect 3004 2892 3068 2956
rect 1825 2748 1889 2752
rect 1825 2692 1829 2748
rect 1829 2692 1885 2748
rect 1885 2692 1889 2748
rect 1825 2688 1889 2692
rect 1905 2748 1969 2752
rect 1905 2692 1909 2748
rect 1909 2692 1965 2748
rect 1965 2692 1969 2748
rect 1905 2688 1969 2692
rect 1985 2748 2049 2752
rect 1985 2692 1989 2748
rect 1989 2692 2045 2748
rect 2045 2692 2049 2748
rect 1985 2688 2049 2692
rect 2065 2748 2129 2752
rect 2065 2692 2069 2748
rect 2069 2692 2125 2748
rect 2125 2692 2129 2748
rect 2065 2688 2129 2692
rect 3572 2748 3636 2752
rect 3572 2692 3576 2748
rect 3576 2692 3632 2748
rect 3632 2692 3636 2748
rect 3572 2688 3636 2692
rect 3652 2748 3716 2752
rect 3652 2692 3656 2748
rect 3656 2692 3712 2748
rect 3712 2692 3716 2748
rect 3652 2688 3716 2692
rect 3732 2748 3796 2752
rect 3732 2692 3736 2748
rect 3736 2692 3792 2748
rect 3792 2692 3796 2748
rect 3732 2688 3796 2692
rect 3812 2748 3876 2752
rect 3812 2692 3816 2748
rect 3816 2692 3872 2748
rect 3872 2692 3876 2748
rect 3812 2688 3876 2692
rect 5319 2748 5383 2752
rect 5319 2692 5323 2748
rect 5323 2692 5379 2748
rect 5379 2692 5383 2748
rect 5319 2688 5383 2692
rect 5399 2748 5463 2752
rect 5399 2692 5403 2748
rect 5403 2692 5459 2748
rect 5459 2692 5463 2748
rect 5399 2688 5463 2692
rect 5479 2748 5543 2752
rect 5479 2692 5483 2748
rect 5483 2692 5539 2748
rect 5539 2692 5543 2748
rect 5479 2688 5543 2692
rect 5559 2748 5623 2752
rect 5559 2692 5563 2748
rect 5563 2692 5619 2748
rect 5619 2692 5623 2748
rect 5559 2688 5623 2692
rect 7066 2748 7130 2752
rect 7066 2692 7070 2748
rect 7070 2692 7126 2748
rect 7126 2692 7130 2748
rect 7066 2688 7130 2692
rect 7146 2748 7210 2752
rect 7146 2692 7150 2748
rect 7150 2692 7206 2748
rect 7206 2692 7210 2748
rect 7146 2688 7210 2692
rect 7226 2748 7290 2752
rect 7226 2692 7230 2748
rect 7230 2692 7286 2748
rect 7286 2692 7290 2748
rect 7226 2688 7290 2692
rect 7306 2748 7370 2752
rect 7306 2692 7310 2748
rect 7310 2692 7366 2748
rect 7366 2692 7370 2748
rect 7306 2688 7370 2692
rect 2485 2204 2549 2208
rect 2485 2148 2489 2204
rect 2489 2148 2545 2204
rect 2545 2148 2549 2204
rect 2485 2144 2549 2148
rect 2565 2204 2629 2208
rect 2565 2148 2569 2204
rect 2569 2148 2625 2204
rect 2625 2148 2629 2204
rect 2565 2144 2629 2148
rect 2645 2204 2709 2208
rect 2645 2148 2649 2204
rect 2649 2148 2705 2204
rect 2705 2148 2709 2204
rect 2645 2144 2709 2148
rect 2725 2204 2789 2208
rect 2725 2148 2729 2204
rect 2729 2148 2785 2204
rect 2785 2148 2789 2204
rect 2725 2144 2789 2148
rect 4232 2204 4296 2208
rect 4232 2148 4236 2204
rect 4236 2148 4292 2204
rect 4292 2148 4296 2204
rect 4232 2144 4296 2148
rect 4312 2204 4376 2208
rect 4312 2148 4316 2204
rect 4316 2148 4372 2204
rect 4372 2148 4376 2204
rect 4312 2144 4376 2148
rect 4392 2204 4456 2208
rect 4392 2148 4396 2204
rect 4396 2148 4452 2204
rect 4452 2148 4456 2204
rect 4392 2144 4456 2148
rect 4472 2204 4536 2208
rect 4472 2148 4476 2204
rect 4476 2148 4532 2204
rect 4532 2148 4536 2204
rect 4472 2144 4536 2148
rect 5979 2204 6043 2208
rect 5979 2148 5983 2204
rect 5983 2148 6039 2204
rect 6039 2148 6043 2204
rect 5979 2144 6043 2148
rect 6059 2204 6123 2208
rect 6059 2148 6063 2204
rect 6063 2148 6119 2204
rect 6119 2148 6123 2204
rect 6059 2144 6123 2148
rect 6139 2204 6203 2208
rect 6139 2148 6143 2204
rect 6143 2148 6199 2204
rect 6199 2148 6203 2204
rect 6139 2144 6203 2148
rect 6219 2204 6283 2208
rect 6219 2148 6223 2204
rect 6223 2148 6279 2204
rect 6279 2148 6283 2204
rect 6219 2144 6283 2148
rect 7726 2204 7790 2208
rect 7726 2148 7730 2204
rect 7730 2148 7786 2204
rect 7786 2148 7790 2204
rect 7726 2144 7790 2148
rect 7806 2204 7870 2208
rect 7806 2148 7810 2204
rect 7810 2148 7866 2204
rect 7866 2148 7870 2204
rect 7806 2144 7870 2148
rect 7886 2204 7950 2208
rect 7886 2148 7890 2204
rect 7890 2148 7946 2204
rect 7946 2148 7950 2204
rect 7886 2144 7950 2148
rect 7966 2204 8030 2208
rect 7966 2148 7970 2204
rect 7970 2148 8026 2204
rect 8026 2148 8030 2204
rect 7966 2144 8030 2148
rect 2268 716 2332 780
<< metal4 >>
rect 1817 8192 2137 8752
rect 1817 8128 1825 8192
rect 1889 8128 1905 8192
rect 1969 8128 1985 8192
rect 2049 8128 2065 8192
rect 2129 8128 2137 8192
rect 1817 7104 2137 8128
rect 1817 7040 1825 7104
rect 1889 7040 1905 7104
rect 1969 7040 1985 7104
rect 2049 7040 2065 7104
rect 2129 7040 2137 7104
rect 1817 6016 2137 7040
rect 2477 8736 2797 8752
rect 2477 8672 2485 8736
rect 2549 8672 2565 8736
rect 2629 8672 2645 8736
rect 2709 8672 2725 8736
rect 2789 8672 2797 8736
rect 2477 7648 2797 8672
rect 2477 7584 2485 7648
rect 2549 7584 2565 7648
rect 2629 7584 2645 7648
rect 2709 7584 2725 7648
rect 2789 7584 2797 7648
rect 2477 6560 2797 7584
rect 2477 6496 2485 6560
rect 2549 6496 2565 6560
rect 2629 6496 2645 6560
rect 2709 6496 2725 6560
rect 2789 6496 2797 6560
rect 2267 6356 2333 6357
rect 2267 6292 2268 6356
rect 2332 6292 2333 6356
rect 2267 6291 2333 6292
rect 1817 5952 1825 6016
rect 1889 5952 1905 6016
rect 1969 5952 1985 6016
rect 2049 5952 2065 6016
rect 2129 5952 2137 6016
rect 1817 4928 2137 5952
rect 1817 4864 1825 4928
rect 1889 4864 1905 4928
rect 1969 4864 1985 4928
rect 2049 4864 2065 4928
rect 2129 4864 2137 4928
rect 1817 3840 2137 4864
rect 1817 3776 1825 3840
rect 1889 3776 1905 3840
rect 1969 3776 1985 3840
rect 2049 3776 2065 3840
rect 2129 3776 2137 3840
rect 1817 2752 2137 3776
rect 1817 2688 1825 2752
rect 1889 2688 1905 2752
rect 1969 2688 1985 2752
rect 2049 2688 2065 2752
rect 2129 2688 2137 2752
rect 1817 2128 2137 2688
rect 2270 781 2330 6291
rect 2477 5472 2797 6496
rect 2477 5408 2485 5472
rect 2549 5408 2565 5472
rect 2629 5408 2645 5472
rect 2709 5408 2725 5472
rect 2789 5408 2797 5472
rect 2477 4384 2797 5408
rect 3564 8192 3884 8752
rect 3564 8128 3572 8192
rect 3636 8128 3652 8192
rect 3716 8128 3732 8192
rect 3796 8128 3812 8192
rect 3876 8128 3884 8192
rect 3564 7104 3884 8128
rect 3564 7040 3572 7104
rect 3636 7040 3652 7104
rect 3716 7040 3732 7104
rect 3796 7040 3812 7104
rect 3876 7040 3884 7104
rect 3564 6016 3884 7040
rect 3564 5952 3572 6016
rect 3636 5952 3652 6016
rect 3716 5952 3732 6016
rect 3796 5952 3812 6016
rect 3876 5952 3884 6016
rect 3003 5132 3069 5133
rect 3003 5068 3004 5132
rect 3068 5068 3069 5132
rect 3003 5067 3069 5068
rect 2477 4320 2485 4384
rect 2549 4320 2565 4384
rect 2629 4320 2645 4384
rect 2709 4320 2725 4384
rect 2789 4320 2797 4384
rect 2477 3296 2797 4320
rect 2477 3232 2485 3296
rect 2549 3232 2565 3296
rect 2629 3232 2645 3296
rect 2709 3232 2725 3296
rect 2789 3232 2797 3296
rect 2477 2208 2797 3232
rect 3006 2957 3066 5067
rect 3564 4928 3884 5952
rect 3564 4864 3572 4928
rect 3636 4864 3652 4928
rect 3716 4864 3732 4928
rect 3796 4864 3812 4928
rect 3876 4864 3884 4928
rect 3564 3840 3884 4864
rect 3564 3776 3572 3840
rect 3636 3776 3652 3840
rect 3716 3776 3732 3840
rect 3796 3776 3812 3840
rect 3876 3776 3884 3840
rect 3003 2956 3069 2957
rect 3003 2892 3004 2956
rect 3068 2892 3069 2956
rect 3003 2891 3069 2892
rect 2477 2144 2485 2208
rect 2549 2144 2565 2208
rect 2629 2144 2645 2208
rect 2709 2144 2725 2208
rect 2789 2144 2797 2208
rect 2477 2128 2797 2144
rect 3564 2752 3884 3776
rect 3564 2688 3572 2752
rect 3636 2688 3652 2752
rect 3716 2688 3732 2752
rect 3796 2688 3812 2752
rect 3876 2688 3884 2752
rect 3564 2128 3884 2688
rect 4224 8736 4544 8752
rect 4224 8672 4232 8736
rect 4296 8672 4312 8736
rect 4376 8672 4392 8736
rect 4456 8672 4472 8736
rect 4536 8672 4544 8736
rect 4224 7648 4544 8672
rect 4224 7584 4232 7648
rect 4296 7584 4312 7648
rect 4376 7584 4392 7648
rect 4456 7584 4472 7648
rect 4536 7584 4544 7648
rect 4224 6560 4544 7584
rect 4224 6496 4232 6560
rect 4296 6496 4312 6560
rect 4376 6496 4392 6560
rect 4456 6496 4472 6560
rect 4536 6496 4544 6560
rect 4224 5472 4544 6496
rect 4224 5408 4232 5472
rect 4296 5408 4312 5472
rect 4376 5408 4392 5472
rect 4456 5408 4472 5472
rect 4536 5408 4544 5472
rect 4224 4384 4544 5408
rect 4224 4320 4232 4384
rect 4296 4320 4312 4384
rect 4376 4320 4392 4384
rect 4456 4320 4472 4384
rect 4536 4320 4544 4384
rect 4224 3296 4544 4320
rect 4224 3232 4232 3296
rect 4296 3232 4312 3296
rect 4376 3232 4392 3296
rect 4456 3232 4472 3296
rect 4536 3232 4544 3296
rect 4224 2208 4544 3232
rect 4224 2144 4232 2208
rect 4296 2144 4312 2208
rect 4376 2144 4392 2208
rect 4456 2144 4472 2208
rect 4536 2144 4544 2208
rect 4224 2128 4544 2144
rect 5311 8192 5631 8752
rect 5311 8128 5319 8192
rect 5383 8128 5399 8192
rect 5463 8128 5479 8192
rect 5543 8128 5559 8192
rect 5623 8128 5631 8192
rect 5311 7104 5631 8128
rect 5311 7040 5319 7104
rect 5383 7040 5399 7104
rect 5463 7040 5479 7104
rect 5543 7040 5559 7104
rect 5623 7040 5631 7104
rect 5311 6016 5631 7040
rect 5311 5952 5319 6016
rect 5383 5952 5399 6016
rect 5463 5952 5479 6016
rect 5543 5952 5559 6016
rect 5623 5952 5631 6016
rect 5311 4928 5631 5952
rect 5311 4864 5319 4928
rect 5383 4864 5399 4928
rect 5463 4864 5479 4928
rect 5543 4864 5559 4928
rect 5623 4864 5631 4928
rect 5311 3840 5631 4864
rect 5311 3776 5319 3840
rect 5383 3776 5399 3840
rect 5463 3776 5479 3840
rect 5543 3776 5559 3840
rect 5623 3776 5631 3840
rect 5311 2752 5631 3776
rect 5311 2688 5319 2752
rect 5383 2688 5399 2752
rect 5463 2688 5479 2752
rect 5543 2688 5559 2752
rect 5623 2688 5631 2752
rect 5311 2128 5631 2688
rect 5971 8736 6291 8752
rect 5971 8672 5979 8736
rect 6043 8672 6059 8736
rect 6123 8672 6139 8736
rect 6203 8672 6219 8736
rect 6283 8672 6291 8736
rect 5971 7648 6291 8672
rect 5971 7584 5979 7648
rect 6043 7584 6059 7648
rect 6123 7584 6139 7648
rect 6203 7584 6219 7648
rect 6283 7584 6291 7648
rect 5971 6560 6291 7584
rect 5971 6496 5979 6560
rect 6043 6496 6059 6560
rect 6123 6496 6139 6560
rect 6203 6496 6219 6560
rect 6283 6496 6291 6560
rect 5971 5472 6291 6496
rect 5971 5408 5979 5472
rect 6043 5408 6059 5472
rect 6123 5408 6139 5472
rect 6203 5408 6219 5472
rect 6283 5408 6291 5472
rect 5971 4384 6291 5408
rect 5971 4320 5979 4384
rect 6043 4320 6059 4384
rect 6123 4320 6139 4384
rect 6203 4320 6219 4384
rect 6283 4320 6291 4384
rect 5971 3296 6291 4320
rect 5971 3232 5979 3296
rect 6043 3232 6059 3296
rect 6123 3232 6139 3296
rect 6203 3232 6219 3296
rect 6283 3232 6291 3296
rect 5971 2208 6291 3232
rect 5971 2144 5979 2208
rect 6043 2144 6059 2208
rect 6123 2144 6139 2208
rect 6203 2144 6219 2208
rect 6283 2144 6291 2208
rect 5971 2128 6291 2144
rect 7058 8192 7378 8752
rect 7058 8128 7066 8192
rect 7130 8128 7146 8192
rect 7210 8128 7226 8192
rect 7290 8128 7306 8192
rect 7370 8128 7378 8192
rect 7058 7104 7378 8128
rect 7058 7040 7066 7104
rect 7130 7040 7146 7104
rect 7210 7040 7226 7104
rect 7290 7040 7306 7104
rect 7370 7040 7378 7104
rect 7058 6016 7378 7040
rect 7058 5952 7066 6016
rect 7130 5952 7146 6016
rect 7210 5952 7226 6016
rect 7290 5952 7306 6016
rect 7370 5952 7378 6016
rect 7058 4928 7378 5952
rect 7058 4864 7066 4928
rect 7130 4864 7146 4928
rect 7210 4864 7226 4928
rect 7290 4864 7306 4928
rect 7370 4864 7378 4928
rect 7058 3840 7378 4864
rect 7058 3776 7066 3840
rect 7130 3776 7146 3840
rect 7210 3776 7226 3840
rect 7290 3776 7306 3840
rect 7370 3776 7378 3840
rect 7058 2752 7378 3776
rect 7058 2688 7066 2752
rect 7130 2688 7146 2752
rect 7210 2688 7226 2752
rect 7290 2688 7306 2752
rect 7370 2688 7378 2752
rect 7058 2128 7378 2688
rect 7718 8736 8038 8752
rect 7718 8672 7726 8736
rect 7790 8672 7806 8736
rect 7870 8672 7886 8736
rect 7950 8672 7966 8736
rect 8030 8672 8038 8736
rect 7718 7648 8038 8672
rect 7718 7584 7726 7648
rect 7790 7584 7806 7648
rect 7870 7584 7886 7648
rect 7950 7584 7966 7648
rect 8030 7584 8038 7648
rect 7718 6560 8038 7584
rect 7718 6496 7726 6560
rect 7790 6496 7806 6560
rect 7870 6496 7886 6560
rect 7950 6496 7966 6560
rect 8030 6496 8038 6560
rect 7718 5472 8038 6496
rect 7718 5408 7726 5472
rect 7790 5408 7806 5472
rect 7870 5408 7886 5472
rect 7950 5408 7966 5472
rect 8030 5408 8038 5472
rect 7718 4384 8038 5408
rect 7718 4320 7726 4384
rect 7790 4320 7806 4384
rect 7870 4320 7886 4384
rect 7950 4320 7966 4384
rect 8030 4320 8038 4384
rect 7718 3296 8038 4320
rect 7718 3232 7726 3296
rect 7790 3232 7806 3296
rect 7870 3232 7886 3296
rect 7950 3232 7966 3296
rect 8030 3232 8038 3296
rect 7718 2208 8038 3232
rect 7718 2144 7726 2208
rect 7790 2144 7806 2208
rect 7870 2144 7886 2208
rect 7950 2144 7966 2208
rect 8030 2144 8038 2208
rect 7718 2128 8038 2144
rect 2267 780 2333 781
rect 2267 716 2268 780
rect 2332 716 2333 780
rect 2267 715 2333 716
use sky130_fd_sc_hd__buf_2  _17_ ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 5152 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1717221846
transform -1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _19_ ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform -1 0 4232 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _20_ ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _21_ ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _22_ ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _23_
timestamp 1717221846
transform -1 0 1840 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1717221846
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _25_
timestamp 1717221846
transform -1 0 4416 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _26_
timestamp 1717221846
transform -1 0 2576 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _27_
timestamp 1717221846
transform -1 0 3680 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1717221846
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _29_
timestamp 1717221846
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _30_
timestamp 1717221846
transform -1 0 2392 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _31_
timestamp 1717221846
transform -1 0 5612 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1717221846
transform -1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _33_
timestamp 1717221846
transform 1 0 1656 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _34_ ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 2484 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _35_
timestamp 1717221846
transform -1 0 2852 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _36_
timestamp 1717221846
transform -1 0 7452 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _37_
timestamp 1717221846
transform -1 0 2484 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _38_
timestamp 1717221846
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _39_
timestamp 1717221846
transform -1 0 7728 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _40_ ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 6532 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _41_
timestamp 1717221846
transform 1 0 5336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _42_
timestamp 1717221846
transform 1 0 7176 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _43_
timestamp 1717221846
transform -1 0 7728 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _44_
timestamp 1717221846
transform -1 0 7636 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _45_
timestamp 1717221846
transform -1 0 2852 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _46_
timestamp 1717221846
transform -1 0 3496 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _47_
timestamp 1717221846
transform 1 0 4508 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _48_ ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1717221846
transform 1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _50_
timestamp 1717221846
transform 1 0 4416 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1717221846
transform -1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _52_
timestamp 1717221846
transform -1 0 4600 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1717221846
transform 1 0 5244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _54_
timestamp 1717221846
transform 1 0 3496 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1717221846
transform 1 0 2576 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _56_ ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 1840 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _57_
timestamp 1717221846
transform 1 0 1840 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _58_
timestamp 1717221846
transform 1 0 4324 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _59_ ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 2392 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _60_ ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 3772 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _61_
timestamp 1717221846
transform -1 0 6808 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _62_
timestamp 1717221846
transform 1 0 5612 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _63_
timestamp 1717221846
transform -1 0 5888 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _64_
timestamp 1717221846
transform 1 0 5888 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _65_
timestamp 1717221846
transform -1 0 7452 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _66_
timestamp 1717221846
transform -1 0 4140 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _67_
timestamp 1717221846
transform 1 0 1840 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform -1 0 6256 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1717221846
transform -1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1717221846
transform 1 0 5244 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1717221846
transform -1 0 5336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_3 ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_7 ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_52
timestamp 1717221846
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69
timestamp 1717221846
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_3
timestamp 1717221846
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_53 ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_57 ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_72
timestamp 1717221846
transform 1 0 7728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3
timestamp 1717221846
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_7
timestamp 1717221846
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_72
timestamp 1717221846
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_3
timestamp 1717221846
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_7
timestamp 1717221846
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1717221846
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_65
timestamp 1717221846
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_15
timestamp 1717221846
transform 1 0 2484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_38
timestamp 1717221846
transform 1 0 4600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_25
timestamp 1717221846
transform 1 0 3404 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_35
timestamp 1717221846
transform 1 0 4324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_61
timestamp 1717221846
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1717221846
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_7
timestamp 1717221846
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_18
timestamp 1717221846
transform 1 0 2760 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1717221846
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 1717221846
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_48
timestamp 1717221846
transform 1 0 5520 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_71
timestamp 1717221846
transform 1 0 7636 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_35 ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 4324 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_43
timestamp 1717221846
transform 1 0 5060 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_69
timestamp 1717221846
transform 1 0 7452 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_33
timestamp 1717221846
transform 1 0 4140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1717221846
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_72
timestamp 1717221846
transform 1 0 7728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_25
timestamp 1717221846
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_37
timestamp 1717221846
transform 1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_15
timestamp 1717221846
transform 1 0 2484 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_29
timestamp 1717221846
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_49 ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1717221846
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1717221846
transform -1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1717221846
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1717221846
transform -1 0 5152 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1717221846
transform -1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1717221846
transform -1 0 7544 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1717221846
transform -1 0 7820 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1717221846
transform -1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1717221846
transform -1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform -1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output2
timestamp 1717221846
transform -1 0 3680 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output3
timestamp 1717221846
transform -1 0 3220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1717221846
transform 1 0 6900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1717221846
transform 1 0 7452 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 1717221846
transform -1 0 3404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output7
timestamp 1717221846
transform -1 0 7820 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 1717221846
transform 1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 1717221846
transform -1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 1717221846
transform 1 0 2852 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1717221846
transform 1 0 4692 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 1717221846
transform -1 0 2484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1717221846
transform -1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1717221846
transform -1 0 4508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1717221846
transform -1 0 2024 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1717221846
transform -1 0 2484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1717221846
transform -1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1717221846
transform 1 0 7452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1717221846
transform -1 0 1932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1717221846
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1717221846
transform 1 0 4232 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1717221846
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1717221846
transform 1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1717221846
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1717221846
transform -1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1717221846
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1717221846
transform -1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1717221846
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1717221846
transform -1 0 8096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1717221846
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1717221846
transform -1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1717221846
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1717221846
transform -1 0 8096 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1717221846
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1717221846
transform -1 0 8096 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1717221846
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1717221846
transform -1 0 8096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1717221846
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1717221846
transform -1 0 8096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1717221846
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1717221846
transform -1 0 8096 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1717221846
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1717221846
transform -1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1717221846
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1717221846
transform -1 0 8096 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1717221846
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1717221846
transform -1 0 8096 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24 ~/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1717221846
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1717221846
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1717221846
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1717221846
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1717221846
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1717221846
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1717221846
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1717221846
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1717221846
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1717221846
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1717221846
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1717221846
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1717221846
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 s 2477 2128 2797 8752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4224 2128 4544 8752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5971 2128 6291 8752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7718 2128 8038 8752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1817 2128 2137 8752 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 3564 2128 3884 8752 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5311 2128 5631 8752 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7058 2128 7378 8752 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 7746 10548 7802 11348 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 ctl0[0]
port 3 nsew signal tristate
flabel metal2 s 2594 10548 2650 11348 0 FreeSans 224 90 0 0 ctl0[1]
port 4 nsew signal tristate
flabel metal3 s 8404 9528 9204 9648 0 FreeSans 480 0 0 0 ctl0[2]
port 5 nsew signal tristate
flabel metal3 s 8404 6128 9204 6248 0 FreeSans 480 0 0 0 ctl0[3]
port 6 nsew signal tristate
flabel metal3 s 8404 2048 9204 2168 0 FreeSans 480 0 0 0 ctl0[4]
port 7 nsew signal tristate
flabel metal2 s 9034 10548 9090 11348 0 FreeSans 224 90 0 0 ctl0[5]
port 8 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 ctl0[6]
port 9 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 ctl0[7]
port 10 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 ctl0[8]
port 11 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 ctl1[0]
port 12 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 ctl1[1]
port 13 nsew signal tristate
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 ctl1[2]
port 14 nsew signal tristate
flabel metal2 s 3882 10548 3938 11348 0 FreeSans 224 90 0 0 ctl1[3]
port 15 nsew signal tristate
flabel metal3 s 8404 688 9204 808 0 FreeSans 480 0 0 0 ctl1[4]
port 16 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 ctl1[5]
port 17 nsew signal tristate
flabel metal2 s 662 10548 718 11348 0 FreeSans 224 90 0 0 ctl1[6]
port 18 nsew signal tristate
flabel metal3 s 8404 7488 9204 7608 0 FreeSans 480 0 0 0 ctl1[7]
port 19 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 ctl1[8]
port 20 nsew signal tristate
flabel metal2 s 5814 10548 5870 11348 0 FreeSans 224 90 0 0 r0_w2_en
port 21 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 r1_w3_en
port 22 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 r2_w0_en
port 23 nsew signal tristate
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 r3_w1_en
port 24 nsew signal tristate
flabel metal3 s 8404 4088 9204 4208 0 FreeSans 480 0 0 0 rst_n
port 25 nsew signal input
rlabel metal1 4600 8704 4600 8704 0 VGND
rlabel metal1 4600 8160 4600 8160 0 VPWR
rlabel metal1 2300 3434 2300 3434 0 _00_
rlabel metal1 2162 2312 2162 2312 0 _01_
rlabel metal1 4646 4216 4646 4216 0 _02_
rlabel metal2 2806 4097 2806 4097 0 _03_
rlabel metal1 1886 7446 1886 7446 0 _04_
rlabel via1 2540 6766 2540 6766 0 _05_
rlabel metal1 3910 2618 3910 2618 0 _06_
rlabel metal1 5888 2414 5888 2414 0 _07_
rlabel metal2 1426 6902 1426 6902 0 _08_
rlabel metal1 1748 4114 1748 4114 0 _09_
rlabel metal1 2162 7888 2162 7888 0 _10_
rlabel metal1 5796 2482 5796 2482 0 _11_
rlabel metal1 4830 7378 4830 7378 0 _12_
rlabel metal1 3036 4454 3036 4454 0 _13_
rlabel metal2 1610 4726 1610 4726 0 _14_
rlabel metal1 4738 4794 4738 4794 0 _15_
rlabel metal1 2898 4590 2898 4590 0 _16_
rlabel metal1 6946 5270 6946 5270 0 clk
rlabel metal1 4692 4998 4692 4998 0 clknet_0_clk
rlabel metal1 2070 2482 2070 2482 0 clknet_1_0__leaf_clk
rlabel metal1 7084 6834 7084 6834 0 clknet_1_1__leaf_clk
rlabel metal3 1717 3468 1717 3468 0 ctl0[0]
rlabel metal2 2714 10064 2714 10064 0 ctl0[1]
rlabel metal2 7130 9095 7130 9095 0 ctl0[2]
rlabel metal1 7912 5882 7912 5882 0 ctl0[3]
rlabel metal3 6555 2380 6555 2380 0 ctl0[4]
rlabel metal1 8326 8602 8326 8602 0 ctl0[5]
rlabel metal2 6486 823 6486 823 0 ctl0[6]
rlabel metal3 820 4828 820 4828 0 ctl0[7]
rlabel metal3 1924 1428 1924 1428 0 ctl0[8]
rlabel metal1 6808 4522 6808 4522 0 ctl1[0]
rlabel metal1 1012 3910 1012 3910 0 ctl1[1]
rlabel metal2 1334 1761 1334 1761 0 ctl1[2]
rlabel metal1 4002 8398 4002 8398 0 ctl1[3]
rlabel metal1 2622 2856 2622 2856 0 ctl1[4]
rlabel metal2 3266 823 3266 823 0 ctl1[5]
rlabel metal1 1518 8296 1518 8296 0 ctl1[6]
rlabel metal1 7912 7718 7912 7718 0 ctl1[7]
rlabel metal3 1096 8908 1096 8908 0 ctl1[8]
rlabel metal1 6571 3434 6571 3434 0 net1
rlabel metal2 3358 4556 3358 4556 0 net10
rlabel metal1 3358 3128 3358 3128 0 net11
rlabel metal1 2300 4590 2300 4590 0 net12
rlabel metal1 1748 4590 1748 4590 0 net13
rlabel metal1 6854 7514 6854 7514 0 net14
rlabel metal1 2714 3026 2714 3026 0 net15
rlabel metal2 1518 5168 1518 5168 0 net16
rlabel metal1 1978 7718 1978 7718 0 net17
rlabel metal1 7498 7922 7498 7922 0 net18
rlabel metal1 1748 7514 1748 7514 0 net19
rlabel metal1 3680 6698 3680 6698 0 net2
rlabel metal1 5198 7242 5198 7242 0 net20
rlabel metal1 4232 2414 4232 2414 0 net21
rlabel metal1 1564 6766 1564 6766 0 net22
rlabel metal1 2116 8058 2116 8058 0 net23
rlabel metal2 3266 2210 3266 2210 0 net24
rlabel metal2 5934 3298 5934 3298 0 net25
rlabel metal1 4278 7310 4278 7310 0 net26
rlabel metal1 6302 7514 6302 7514 0 net27
rlabel metal1 4278 5882 4278 5882 0 net28
rlabel metal2 2254 6154 2254 6154 0 net29
rlabel metal2 3082 7548 3082 7548 0 net3
rlabel metal1 7176 5338 7176 5338 0 net30
rlabel metal1 5704 3434 5704 3434 0 net31
rlabel metal2 5934 6392 5934 6392 0 net32
rlabel metal2 6394 4454 6394 4454 0 net33
rlabel metal2 6854 8262 6854 8262 0 net4
rlabel metal1 7682 5678 7682 5678 0 net5
rlabel metal2 6578 5236 6578 5236 0 net6
rlabel metal1 7682 4250 7682 4250 0 net7
rlabel metal1 6992 2414 6992 2414 0 net8
rlabel metal1 1932 5270 1932 5270 0 net9
rlabel metal2 3634 3162 3634 3162 0 phase\[0\]
rlabel metal1 3634 2448 3634 2448 0 phase\[1\]
rlabel metal1 6670 5134 6670 5134 0 phase\[2\]
rlabel metal1 6486 2312 6486 2312 0 phase\[3\]
rlabel metal1 6210 8602 6210 8602 0 r0_w2_en
rlabel metal2 5198 959 5198 959 0 r1_w3_en
rlabel metal3 820 6868 820 6868 0 r2_w0_en
rlabel metal2 2898 9401 2898 9401 0 r3_w1_en
rlabel metal1 7958 5202 7958 5202 0 rst_n
rlabel metal2 3082 5406 3082 5406 0 step\[0\]
rlabel metal1 2346 7854 2346 7854 0 step\[1\]
rlabel metal1 6762 6222 6762 6222 0 step\[2\]
rlabel metal2 5290 3196 5290 3196 0 step\[3\]
rlabel metal1 6854 6358 6854 6358 0 step\[4\]
rlabel viali 2622 7852 2622 7852 0 step\[5\]
rlabel metal1 2576 6698 2576 6698 0 step\[6\]
rlabel metal1 4094 5168 4094 5168 0 step\[7\]
<< properties >>
string FIXED_BBOX 0 0 9204 11348
<< end >>
