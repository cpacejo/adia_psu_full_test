VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_adia_psu_full_test
  CLASS BLOCK ;
  FOREIGN tt_um_adia_psu_full_test ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.912600 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.310500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.310500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.310500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.310500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.310500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.310500 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.310500 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.054499 ;
    ANTENNADIFFAREA 114.046097 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.054499 ;
    ANTENNADIFFAREA 114.046097 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.054499 ;
    ANTENNADIFFAREA 114.046097 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.054499 ;
    ANTENNADIFFAREA 114.046097 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.054499 ;
    ANTENNADIFFAREA 114.046097 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.054499 ;
    ANTENNADIFFAREA 114.046097 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.054499 ;
    ANTENNADIFFAREA 114.046097 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.054499 ;
    ANTENNADIFFAREA 114.046097 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.063000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 25.395300 ;
    ANTENNADIFFAREA 72.564751 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.063000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.063000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.310500 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.310500 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.310500 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 8.415 207.415 8.585 207.605 ;
        RECT 12.095 207.415 12.265 207.605 ;
        RECT 12.555 207.415 12.725 207.605 ;
        RECT 15.325 207.460 15.485 207.570 ;
        RECT 18.535 207.415 18.705 207.605 ;
        RECT 20.835 207.435 21.005 207.605 ;
        RECT 21.765 207.460 21.925 207.570 ;
        RECT 20.835 207.415 20.985 207.435 ;
        RECT 24.975 207.415 25.145 207.605 ;
        RECT 25.435 207.415 25.605 207.605 ;
        RECT 30.495 207.435 30.665 207.605 ;
        RECT 30.495 207.415 30.645 207.435 ;
        RECT 30.955 207.415 31.125 207.605 ;
        RECT 33.710 207.465 33.830 207.575 ;
        RECT 34.635 207.415 34.805 207.605 ;
        RECT 37.395 207.415 37.565 207.605 ;
        RECT 41.535 207.415 41.705 207.605 ;
        RECT 42.915 207.415 43.085 207.605 ;
        RECT 8.275 206.605 9.645 207.415 ;
        RECT 9.665 206.735 12.405 207.415 ;
        RECT 12.415 206.735 15.155 207.415 ;
        RECT 16.105 206.735 18.845 207.415 ;
        RECT 19.055 206.595 20.985 207.415 ;
        RECT 19.055 206.505 20.005 206.595 ;
        RECT 21.165 206.545 21.595 207.330 ;
        RECT 22.545 206.735 25.285 207.415 ;
        RECT 25.295 206.505 28.505 207.415 ;
        RECT 28.715 206.595 30.645 207.415 ;
        RECT 30.815 206.605 33.565 207.415 ;
        RECT 28.715 206.505 29.665 206.595 ;
        RECT 34.045 206.545 34.475 207.330 ;
        RECT 34.495 206.735 37.235 207.415 ;
        RECT 37.255 206.735 39.085 207.415 ;
        RECT 39.105 206.735 41.845 207.415 ;
        RECT 37.740 206.505 39.085 206.735 ;
        RECT 41.855 206.605 43.225 207.415 ;
      LAYER nwell ;
        RECT 8.080 203.385 43.420 206.215 ;
      LAYER pwell ;
        RECT 8.275 202.185 9.645 202.995 ;
        RECT 9.665 202.185 12.405 202.865 ;
        RECT 12.415 202.185 13.785 202.965 ;
        RECT 13.795 202.185 17.005 203.095 ;
        RECT 17.025 202.185 19.765 202.865 ;
        RECT 19.775 202.185 21.145 202.995 ;
        RECT 21.165 202.270 21.595 203.055 ;
        RECT 21.710 202.865 22.630 203.095 ;
        RECT 21.710 202.185 25.175 202.865 ;
        RECT 25.295 202.185 27.125 202.995 ;
        RECT 27.175 202.865 28.515 203.095 ;
        RECT 31.345 202.865 32.275 203.085 ;
        RECT 27.175 202.185 36.785 202.865 ;
        RECT 36.795 202.185 40.005 203.095 ;
        RECT 40.500 202.865 41.845 203.095 ;
        RECT 40.015 202.185 41.845 202.865 ;
        RECT 41.855 202.185 43.225 202.995 ;
        RECT 8.415 201.975 8.585 202.185 ;
        RECT 9.795 201.975 9.965 202.165 ;
        RECT 11.175 201.975 11.345 202.165 ;
        RECT 12.095 201.995 12.265 202.185 ;
        RECT 13.475 201.995 13.645 202.185 ;
        RECT 16.695 201.995 16.865 202.185 ;
        RECT 19.455 201.995 19.625 202.185 ;
        RECT 19.915 201.995 20.085 202.185 ;
        RECT 23.135 201.975 23.305 202.165 ;
        RECT 23.595 201.975 23.765 202.165 ;
        RECT 24.975 201.975 25.145 202.185 ;
        RECT 25.435 201.995 25.605 202.185 ;
        RECT 29.575 201.975 29.745 202.165 ;
        RECT 30.035 201.975 30.205 202.165 ;
        RECT 33.710 202.025 33.830 202.135 ;
        RECT 36.475 201.995 36.645 202.185 ;
        RECT 37.855 201.975 38.025 202.165 ;
        RECT 39.695 201.995 39.865 202.185 ;
        RECT 40.155 201.995 40.325 202.185 ;
        RECT 41.075 201.975 41.245 202.165 ;
        RECT 41.530 202.025 41.650 202.135 ;
        RECT 42.915 201.975 43.085 202.185 ;
        RECT 8.275 201.165 9.645 201.975 ;
        RECT 9.655 201.195 11.025 201.975 ;
        RECT 11.045 201.065 13.775 201.975 ;
        RECT 13.835 201.295 23.445 201.975 ;
        RECT 13.835 201.065 15.175 201.295 ;
        RECT 18.005 201.075 18.935 201.295 ;
        RECT 23.455 201.165 24.825 201.975 ;
        RECT 24.835 201.195 26.205 201.975 ;
        RECT 26.310 201.295 29.775 201.975 ;
        RECT 30.005 201.295 33.470 201.975 ;
        RECT 26.310 201.065 27.230 201.295 ;
        RECT 32.550 201.065 33.470 201.295 ;
        RECT 34.045 201.105 34.475 201.890 ;
        RECT 34.590 201.295 38.055 201.975 ;
        RECT 34.590 201.065 35.510 201.295 ;
        RECT 38.175 201.065 41.385 201.975 ;
        RECT 41.855 201.165 43.225 201.975 ;
      LAYER nwell ;
        RECT 8.080 197.945 43.420 200.775 ;
      LAYER pwell ;
        RECT 8.275 196.745 9.645 197.555 ;
        RECT 9.655 196.745 12.395 197.425 ;
        RECT 12.425 196.745 15.165 197.425 ;
        RECT 15.175 196.745 18.385 197.655 ;
        RECT 18.405 196.745 21.145 197.425 ;
        RECT 21.165 196.830 21.595 197.615 ;
        RECT 21.625 196.745 24.355 197.655 ;
        RECT 24.375 196.745 28.045 197.555 ;
        RECT 28.975 196.745 30.345 197.525 ;
        RECT 30.395 197.425 31.735 197.655 ;
        RECT 34.565 197.425 35.495 197.645 ;
        RECT 30.395 196.745 40.005 197.425 ;
        RECT 40.015 196.745 41.845 197.555 ;
        RECT 41.855 196.745 43.225 197.555 ;
        RECT 8.415 196.535 8.585 196.745 ;
        RECT 9.795 196.555 9.965 196.745 ;
        RECT 11.635 196.555 11.805 196.725 ;
        RECT 11.635 196.535 11.785 196.555 ;
        RECT 12.095 196.535 12.265 196.725 ;
        RECT 14.855 196.555 15.025 196.745 ;
        RECT 15.315 196.555 15.485 196.745 ;
        RECT 20.835 196.555 21.005 196.745 ;
        RECT 21.755 196.535 21.925 196.745 ;
        RECT 24.515 196.555 24.685 196.745 ;
        RECT 28.205 196.590 28.365 196.700 ;
        RECT 30.035 196.555 30.205 196.745 ;
        RECT 31.415 196.535 31.585 196.725 ;
        RECT 34.635 196.535 34.805 196.725 ;
        RECT 39.695 196.555 39.865 196.745 ;
        RECT 40.155 196.555 40.325 196.745 ;
        RECT 40.615 196.535 40.785 196.725 ;
        RECT 41.085 196.580 41.245 196.690 ;
        RECT 42.915 196.535 43.085 196.745 ;
        RECT 8.275 195.725 9.645 196.535 ;
        RECT 9.855 195.715 11.785 196.535 ;
        RECT 11.955 195.855 21.235 196.535 ;
        RECT 21.615 195.855 31.225 196.535 ;
        RECT 31.275 195.855 34.015 196.535 ;
        RECT 9.855 195.625 10.805 195.715 ;
        RECT 13.315 195.635 14.235 195.855 ;
        RECT 18.900 195.735 21.235 195.855 ;
        RECT 20.315 195.625 21.235 195.735 ;
        RECT 26.125 195.635 27.055 195.855 ;
        RECT 29.885 195.625 31.225 195.855 ;
        RECT 34.045 195.665 34.475 196.450 ;
        RECT 34.495 195.625 37.705 196.535 ;
        RECT 37.715 195.625 40.925 196.535 ;
        RECT 41.855 195.725 43.225 196.535 ;
      LAYER nwell ;
        RECT 8.080 192.505 43.420 195.335 ;
      LAYER pwell ;
        RECT 8.275 191.305 9.645 192.115 ;
        RECT 9.655 191.305 11.485 192.115 ;
        RECT 11.955 191.305 15.165 192.215 ;
        RECT 15.175 191.305 16.545 192.085 ;
        RECT 17.015 191.305 20.225 192.215 ;
        RECT 21.165 191.390 21.595 192.175 ;
        RECT 24.930 191.985 25.850 192.215 ;
        RECT 29.000 191.985 30.345 192.215 ;
        RECT 35.325 191.985 36.255 192.205 ;
        RECT 39.085 191.985 40.005 192.215 ;
        RECT 40.500 191.985 41.845 192.215 ;
        RECT 22.085 191.305 24.825 191.985 ;
        RECT 24.930 191.305 28.395 191.985 ;
        RECT 28.515 191.305 30.345 191.985 ;
        RECT 30.815 191.305 40.005 191.985 ;
        RECT 40.015 191.305 41.845 191.985 ;
        RECT 41.855 191.305 43.225 192.115 ;
        RECT 8.415 191.095 8.585 191.305 ;
        RECT 9.795 191.115 9.965 191.305 ;
        RECT 11.630 191.145 11.750 191.255 ;
        RECT 12.095 191.095 12.265 191.285 ;
        RECT 12.555 191.095 12.725 191.285 ;
        RECT 14.855 191.115 15.025 191.305 ;
        RECT 16.235 191.115 16.405 191.305 ;
        RECT 16.695 191.255 16.865 191.285 ;
        RECT 16.690 191.145 16.865 191.255 ;
        RECT 16.695 191.095 16.865 191.145 ;
        RECT 17.155 191.095 17.325 191.285 ;
        RECT 19.915 191.255 20.085 191.305 ;
        RECT 19.910 191.145 20.085 191.255 ;
        RECT 20.385 191.150 20.545 191.260 ;
        RECT 19.915 191.115 20.085 191.145 ;
        RECT 20.650 191.095 20.820 191.285 ;
        RECT 24.515 191.255 24.685 191.305 ;
        RECT 21.750 191.145 21.870 191.255 ;
        RECT 24.510 191.145 24.685 191.255 ;
        RECT 24.515 191.115 24.685 191.145 ;
        RECT 28.195 191.115 28.365 191.305 ;
        RECT 28.655 191.115 28.825 191.305 ;
        RECT 30.490 191.145 30.610 191.255 ;
        RECT 30.955 191.115 31.125 191.305 ;
        RECT 33.715 191.095 33.885 191.285 ;
        RECT 36.015 191.095 36.185 191.285 ;
        RECT 36.470 191.145 36.590 191.255 ;
        RECT 40.155 191.095 40.325 191.305 ;
        RECT 41.525 191.095 41.695 191.285 ;
        RECT 42.915 191.095 43.085 191.305 ;
        RECT 8.275 190.285 9.645 191.095 ;
        RECT 9.665 190.415 12.405 191.095 ;
        RECT 12.415 190.315 13.785 191.095 ;
        RECT 13.795 190.185 17.005 191.095 ;
        RECT 17.015 190.415 19.755 191.095 ;
        RECT 20.235 190.415 24.135 191.095 ;
        RECT 24.920 190.415 34.025 191.095 ;
        RECT 20.235 190.185 21.165 190.415 ;
        RECT 34.045 190.225 34.475 191.010 ;
        RECT 34.495 190.415 36.325 191.095 ;
        RECT 36.890 190.415 40.355 191.095 ;
        RECT 34.495 190.185 35.840 190.415 ;
        RECT 36.890 190.185 37.810 190.415 ;
        RECT 40.475 190.315 41.845 191.095 ;
        RECT 41.855 190.285 43.225 191.095 ;
      LAYER nwell ;
        RECT 8.080 187.065 43.420 189.895 ;
        RECT 59.980 188.235 62.290 190.815 ;
      LAYER pwell ;
        RECT 8.275 185.865 9.645 186.675 ;
        RECT 9.665 185.865 12.405 186.545 ;
        RECT 12.425 185.865 15.165 186.545 ;
        RECT 15.635 185.865 17.005 186.645 ;
        RECT 17.015 186.545 17.945 186.775 ;
        RECT 17.015 185.865 20.915 186.545 ;
        RECT 21.165 185.950 21.595 186.735 ;
        RECT 24.815 186.545 25.745 186.775 ;
        RECT 38.270 186.545 39.190 186.775 ;
        RECT 21.845 185.865 25.745 186.545 ;
        RECT 26.215 185.865 28.955 186.545 ;
        RECT 28.975 185.865 38.080 186.545 ;
        RECT 38.270 185.865 41.735 186.545 ;
        RECT 41.855 185.865 43.225 186.675 ;
      LAYER nwell ;
        RECT 58.320 186.630 62.290 188.235 ;
        RECT 59.980 186.625 62.290 186.630 ;
      LAYER pwell ;
        RECT 8.415 185.655 8.585 185.865 ;
        RECT 9.795 185.655 9.965 185.845 ;
        RECT 11.630 185.705 11.750 185.815 ;
        RECT 12.095 185.675 12.265 185.865 ;
        RECT 14.395 185.655 14.565 185.845 ;
        RECT 14.855 185.655 15.025 185.865 ;
        RECT 15.310 185.705 15.430 185.815 ;
        RECT 16.695 185.675 16.865 185.865 ;
        RECT 17.430 185.675 17.600 185.865 ;
        RECT 24.515 185.655 24.685 185.845 ;
        RECT 25.160 185.675 25.330 185.865 ;
        RECT 25.890 185.705 26.010 185.815 ;
        RECT 26.355 185.675 26.525 185.865 ;
        RECT 29.115 185.675 29.285 185.865 ;
        RECT 33.710 185.705 33.830 185.815 ;
        RECT 37.855 185.655 38.025 185.845 ;
        RECT 38.310 185.705 38.430 185.815 ;
        RECT 38.775 185.655 38.945 185.845 ;
        RECT 41.535 185.675 41.705 185.865 ;
        RECT 42.915 185.655 43.085 185.865 ;
        RECT 8.275 184.845 9.645 185.655 ;
        RECT 9.655 184.845 11.485 185.655 ;
        RECT 11.965 184.745 14.695 185.655 ;
        RECT 14.715 184.975 23.995 185.655 ;
        RECT 24.375 184.975 33.565 185.655 ;
        RECT 16.075 184.755 16.995 184.975 ;
        RECT 21.660 184.855 23.995 184.975 ;
        RECT 23.075 184.745 23.995 184.855 ;
        RECT 28.885 184.755 29.815 184.975 ;
        RECT 32.645 184.745 33.565 184.975 ;
        RECT 34.045 184.785 34.475 185.570 ;
        RECT 34.590 184.975 38.055 185.655 ;
        RECT 34.590 184.745 35.510 184.975 ;
        RECT 38.635 184.745 41.845 185.655 ;
        RECT 41.855 184.845 43.225 185.655 ;
        RECT 58.720 185.430 59.650 186.340 ;
        RECT 58.720 185.410 58.825 185.430 ;
        RECT 58.655 185.240 58.825 185.410 ;
      LAYER nwell ;
        RECT 8.080 181.625 43.420 184.455 ;
      LAYER pwell ;
        RECT 60.090 184.035 62.200 186.555 ;
        RECT 8.275 180.425 9.645 181.235 ;
        RECT 9.655 180.425 11.485 181.235 ;
        RECT 16.465 181.105 17.395 181.325 ;
        RECT 20.225 181.105 21.145 181.335 ;
        RECT 11.955 180.425 21.145 181.105 ;
        RECT 21.165 180.510 21.595 181.295 ;
        RECT 21.615 180.425 22.985 181.205 ;
        RECT 22.995 181.105 23.915 181.335 ;
        RECT 26.745 181.105 27.675 181.325 ;
        RECT 36.705 181.105 37.635 181.325 ;
        RECT 40.465 181.105 41.385 181.335 ;
        RECT 22.995 180.425 32.185 181.105 ;
        RECT 32.195 180.425 41.385 181.105 ;
        RECT 41.855 180.425 43.225 181.235 ;
        RECT 8.415 180.215 8.585 180.425 ;
        RECT 9.795 180.375 9.965 180.425 ;
        RECT 9.790 180.265 9.965 180.375 ;
        RECT 11.630 180.265 11.750 180.375 ;
        RECT 9.795 180.235 9.965 180.265 ;
        RECT 12.095 180.235 12.265 180.425 ;
        RECT 12.555 180.215 12.725 180.405 ;
        RECT 15.315 180.215 15.485 180.405 ;
        RECT 21.755 180.235 21.925 180.425 ;
        RECT 24.515 180.215 24.685 180.405 ;
        RECT 25.250 180.215 25.420 180.405 ;
        RECT 29.115 180.215 29.285 180.405 ;
        RECT 31.875 180.235 32.045 180.425 ;
        RECT 32.335 180.235 32.505 180.425 ;
        RECT 32.795 180.215 32.965 180.405 ;
        RECT 34.645 180.260 34.805 180.370 ;
        RECT 35.555 180.215 35.725 180.405 ;
        RECT 41.075 180.215 41.245 180.405 ;
        RECT 41.530 180.265 41.650 180.375 ;
        RECT 42.915 180.215 43.085 180.425 ;
        RECT 8.275 179.405 9.645 180.215 ;
        RECT 10.125 179.535 12.865 180.215 ;
        RECT 12.885 179.305 15.615 180.215 ;
        RECT 15.720 179.535 24.825 180.215 ;
        RECT 24.835 179.535 28.735 180.215 ;
        RECT 29.085 179.535 32.550 180.215 ;
        RECT 24.835 179.305 25.765 179.535 ;
        RECT 31.630 179.305 32.550 179.535 ;
        RECT 32.655 179.405 34.025 180.215 ;
        RECT 34.045 179.345 34.475 180.130 ;
        RECT 35.415 179.305 38.165 180.215 ;
        RECT 38.175 179.305 41.385 180.215 ;
        RECT 41.855 179.405 43.225 180.215 ;
      LAYER nwell ;
        RECT 8.080 176.185 43.420 179.015 ;
      LAYER pwell ;
        RECT 8.275 174.985 9.645 175.795 ;
        RECT 9.655 174.985 11.485 175.795 ;
        RECT 16.465 175.665 17.395 175.885 ;
        RECT 20.225 175.665 21.145 175.895 ;
        RECT 11.955 174.985 21.145 175.665 ;
        RECT 21.165 175.070 21.595 175.855 ;
        RECT 21.815 175.805 22.765 175.895 ;
        RECT 21.815 174.985 23.745 175.805 ;
        RECT 23.915 174.985 26.655 175.665 ;
        RECT 26.685 174.985 29.425 175.665 ;
        RECT 29.435 174.985 32.185 175.895 ;
        RECT 32.195 174.985 34.025 175.795 ;
        RECT 34.045 175.070 34.475 175.855 ;
        RECT 34.495 174.985 37.235 175.665 ;
        RECT 37.255 174.985 39.995 175.665 ;
        RECT 40.015 174.985 41.845 175.795 ;
        RECT 41.855 174.985 43.225 175.795 ;
        RECT 8.415 174.795 8.585 174.985 ;
        RECT 9.795 174.795 9.965 174.985 ;
        RECT 11.630 174.825 11.750 174.935 ;
        RECT 12.095 174.795 12.265 174.985 ;
        RECT 23.595 174.965 23.745 174.985 ;
        RECT 23.595 174.795 23.765 174.965 ;
        RECT 24.055 174.795 24.225 174.985 ;
        RECT 29.115 174.795 29.285 174.985 ;
        RECT 29.575 174.795 29.745 174.985 ;
        RECT 32.335 174.795 32.505 174.985 ;
        RECT 34.635 174.795 34.805 174.985 ;
        RECT 37.395 174.795 37.565 174.985 ;
        RECT 40.155 174.795 40.325 174.985 ;
        RECT 42.915 174.795 43.085 174.985 ;
      LAYER nwell ;
        RECT 58.775 158.765 61.085 161.345 ;
        RECT 57.115 157.160 61.085 158.765 ;
        RECT 58.775 157.155 61.085 157.160 ;
      LAYER pwell ;
        RECT 57.515 155.960 58.445 156.870 ;
        RECT 57.515 155.940 57.620 155.960 ;
        RECT 57.450 155.770 57.620 155.940 ;
        RECT 58.885 154.565 60.995 157.085 ;
      LAYER nwell ;
        RECT 58.610 128.935 60.920 131.515 ;
        RECT 56.950 127.330 60.920 128.935 ;
        RECT 58.610 127.325 60.920 127.330 ;
      LAYER pwell ;
        RECT 57.350 126.130 58.280 127.040 ;
        RECT 57.350 126.110 57.455 126.130 ;
        RECT 57.285 125.940 57.455 126.110 ;
        RECT 58.720 124.735 60.830 127.255 ;
      LAYER nwell ;
        RECT 19.720 102.330 22.030 104.910 ;
        RECT 18.060 100.725 22.030 102.330 ;
      LAYER pwell ;
        RECT 34.780 101.140 37.300 103.250 ;
        RECT 39.820 101.130 42.340 103.240 ;
        RECT 44.780 101.120 47.300 103.230 ;
      LAYER nwell ;
        RECT 19.720 100.720 22.030 100.725 ;
      LAYER pwell ;
        RECT 18.460 99.525 19.390 100.435 ;
        RECT 18.460 99.505 18.565 99.525 ;
        RECT 18.395 99.335 18.565 99.505 ;
        RECT 19.830 98.130 21.940 100.650 ;
      LAYER nwell ;
        RECT 59.070 98.075 61.380 100.655 ;
        RECT 57.410 96.470 61.380 98.075 ;
        RECT 59.070 96.465 61.380 96.470 ;
      LAYER pwell ;
        RECT 57.810 95.270 58.740 96.180 ;
        RECT 57.810 95.250 57.915 95.270 ;
        RECT 57.745 95.080 57.915 95.250 ;
        RECT 59.180 93.875 61.290 96.395 ;
      LAYER nwell ;
        RECT 19.870 91.260 22.180 93.840 ;
        RECT 18.210 89.655 22.180 91.260 ;
        RECT 19.870 89.650 22.180 89.655 ;
      LAYER pwell ;
        RECT 18.610 88.455 19.540 89.365 ;
        RECT 18.610 88.435 18.715 88.455 ;
        RECT 18.545 88.265 18.715 88.435 ;
        RECT 19.980 87.060 22.090 89.580 ;
      LAYER nwell ;
        RECT 19.820 80.130 22.130 82.710 ;
        RECT 18.160 78.525 22.130 80.130 ;
        RECT 28.585 79.430 31.775 79.910 ;
        RECT 19.820 78.520 22.130 78.525 ;
      LAYER pwell ;
        RECT 18.560 77.325 19.490 78.235 ;
        RECT 18.560 77.305 18.665 77.325 ;
        RECT 18.495 77.135 18.665 77.305 ;
        RECT 19.930 75.930 22.040 78.450 ;
      LAYER nwell ;
        RECT 26.850 77.825 31.775 79.430 ;
        RECT 36.135 79.375 39.325 79.855 ;
        RECT 43.130 79.375 46.320 79.855 ;
        RECT 28.585 77.800 31.775 77.825 ;
        RECT 34.400 77.770 39.325 79.375 ;
        RECT 41.395 77.770 46.320 79.375 ;
        RECT 36.135 77.745 39.325 77.770 ;
        RECT 43.130 77.745 46.320 77.770 ;
      LAYER pwell ;
        RECT 27.250 76.625 28.180 77.535 ;
        RECT 27.250 76.605 27.355 76.625 ;
        RECT 27.185 76.435 27.355 76.605 ;
        RECT 34.800 76.570 35.730 77.480 ;
        RECT 41.795 76.570 42.725 77.480 ;
        RECT 34.800 76.550 34.905 76.570 ;
        RECT 41.795 76.550 41.900 76.570 ;
        RECT 34.735 76.380 34.905 76.550 ;
        RECT 41.730 76.380 41.900 76.550 ;
      LAYER nwell ;
        RECT 58.570 68.310 60.880 70.890 ;
        RECT 56.910 66.705 60.880 68.310 ;
        RECT 58.570 66.700 60.880 66.705 ;
      LAYER pwell ;
        RECT 57.310 65.505 58.240 66.415 ;
        RECT 57.310 65.485 57.415 65.505 ;
        RECT 57.245 65.315 57.415 65.485 ;
        RECT 58.680 64.110 60.790 66.630 ;
      LAYER nwell ;
        RECT 58.440 38.815 60.750 41.395 ;
        RECT 56.780 37.210 60.750 38.815 ;
        RECT 58.440 37.205 60.750 37.210 ;
      LAYER pwell ;
        RECT 57.180 36.010 58.110 36.920 ;
        RECT 57.180 35.990 57.285 36.010 ;
        RECT 57.115 35.820 57.285 35.990 ;
        RECT 58.550 34.615 60.660 37.135 ;
      LAYER nwell ;
        RECT 59.470 7.100 61.780 9.680 ;
        RECT 57.810 5.495 61.780 7.100 ;
        RECT 59.470 5.490 61.780 5.495 ;
      LAYER pwell ;
        RECT 58.210 4.295 59.140 5.205 ;
        RECT 58.210 4.275 58.315 4.295 ;
        RECT 58.145 4.105 58.315 4.275 ;
        RECT 59.580 2.900 61.690 5.420 ;
      LAYER li1 ;
        RECT 8.270 207.435 43.230 207.605 ;
        RECT 8.355 206.685 9.565 207.435 ;
        RECT 9.795 206.955 10.075 207.435 ;
        RECT 10.245 206.785 10.505 207.175 ;
        RECT 10.680 206.955 10.935 207.435 ;
        RECT 11.105 206.785 11.400 207.175 ;
        RECT 11.580 206.955 11.855 207.435 ;
        RECT 12.025 206.935 12.325 207.265 ;
        RECT 8.355 206.145 8.875 206.685 ;
        RECT 9.750 206.615 11.400 206.785 ;
        RECT 9.045 205.975 9.565 206.515 ;
        RECT 8.355 204.885 9.565 205.975 ;
        RECT 9.750 206.105 10.155 206.615 ;
        RECT 10.325 206.275 11.465 206.445 ;
        RECT 9.750 205.935 10.505 206.105 ;
        RECT 9.790 204.885 10.075 205.755 ;
        RECT 10.245 205.685 10.505 205.935 ;
        RECT 11.295 206.025 11.465 206.275 ;
        RECT 11.635 206.195 11.985 206.765 ;
        RECT 12.155 206.025 12.325 206.935 ;
        RECT 11.295 205.855 12.325 206.025 ;
        RECT 10.245 205.515 11.365 205.685 ;
        RECT 10.245 205.055 10.505 205.515 ;
        RECT 10.680 204.885 10.935 205.345 ;
        RECT 11.105 205.055 11.365 205.515 ;
        RECT 11.535 204.885 11.845 205.685 ;
        RECT 12.015 205.055 12.325 205.855 ;
        RECT 12.495 206.935 12.795 207.265 ;
        RECT 12.965 206.955 13.240 207.435 ;
        RECT 12.495 206.025 12.665 206.935 ;
        RECT 13.420 206.785 13.715 207.175 ;
        RECT 13.885 206.955 14.140 207.435 ;
        RECT 14.315 206.785 14.575 207.175 ;
        RECT 14.745 206.955 15.025 207.435 ;
        RECT 16.235 206.955 16.515 207.435 ;
        RECT 16.685 206.785 16.945 207.175 ;
        RECT 17.120 206.955 17.375 207.435 ;
        RECT 17.545 206.785 17.840 207.175 ;
        RECT 18.020 206.955 18.295 207.435 ;
        RECT 18.465 206.935 18.765 207.265 ;
        RECT 12.835 206.195 13.185 206.765 ;
        RECT 13.420 206.615 15.070 206.785 ;
        RECT 13.355 206.275 14.495 206.445 ;
        RECT 13.355 206.025 13.525 206.275 ;
        RECT 14.665 206.105 15.070 206.615 ;
        RECT 12.495 205.855 13.525 206.025 ;
        RECT 14.315 205.935 15.070 206.105 ;
        RECT 16.190 206.615 17.840 206.785 ;
        RECT 16.190 206.105 16.595 206.615 ;
        RECT 16.765 206.275 17.905 206.445 ;
        RECT 16.190 205.935 16.945 206.105 ;
        RECT 12.495 205.055 12.805 205.855 ;
        RECT 14.315 205.685 14.575 205.935 ;
        RECT 12.975 204.885 13.285 205.685 ;
        RECT 13.455 205.515 14.575 205.685 ;
        RECT 13.455 205.055 13.715 205.515 ;
        RECT 13.885 204.885 14.140 205.345 ;
        RECT 14.315 205.055 14.575 205.515 ;
        RECT 14.745 204.885 15.030 205.755 ;
        RECT 16.230 204.885 16.515 205.755 ;
        RECT 16.685 205.685 16.945 205.935 ;
        RECT 17.735 206.025 17.905 206.275 ;
        RECT 18.075 206.195 18.425 206.765 ;
        RECT 18.595 206.025 18.765 206.935 ;
        RECT 17.735 205.855 18.765 206.025 ;
        RECT 16.685 205.515 17.805 205.685 ;
        RECT 16.685 205.055 16.945 205.515 ;
        RECT 17.120 204.885 17.375 205.345 ;
        RECT 17.545 205.055 17.805 205.515 ;
        RECT 17.975 204.885 18.285 205.685 ;
        RECT 18.455 205.055 18.765 205.855 ;
        RECT 18.935 206.975 19.495 207.265 ;
        RECT 19.665 206.975 19.915 207.435 ;
        RECT 18.935 205.605 19.185 206.975 ;
        RECT 20.535 206.805 20.865 207.165 ;
        RECT 19.475 206.615 20.865 206.805 ;
        RECT 21.235 206.710 21.525 207.435 ;
        RECT 22.675 206.955 22.955 207.435 ;
        RECT 23.125 206.785 23.385 207.175 ;
        RECT 23.560 206.955 23.815 207.435 ;
        RECT 23.985 206.785 24.280 207.175 ;
        RECT 24.460 206.955 24.735 207.435 ;
        RECT 24.905 206.935 25.205 207.265 ;
        RECT 22.630 206.615 24.280 206.785 ;
        RECT 19.475 206.525 19.645 206.615 ;
        RECT 19.355 206.195 19.645 206.525 ;
        RECT 19.815 206.195 20.155 206.445 ;
        RECT 20.375 206.195 21.050 206.445 ;
        RECT 19.475 205.945 19.645 206.195 ;
        RECT 19.475 205.775 20.415 205.945 ;
        RECT 20.785 205.835 21.050 206.195 ;
        RECT 22.630 206.105 23.035 206.615 ;
        RECT 23.205 206.275 24.345 206.445 ;
        RECT 18.935 205.055 19.395 205.605 ;
        RECT 19.585 204.885 19.915 205.605 ;
        RECT 20.115 205.225 20.415 205.775 ;
        RECT 20.585 204.885 20.865 205.555 ;
        RECT 21.235 204.885 21.525 206.050 ;
        RECT 22.630 205.935 23.385 206.105 ;
        RECT 22.670 204.885 22.955 205.755 ;
        RECT 23.125 205.685 23.385 205.935 ;
        RECT 24.175 206.025 24.345 206.275 ;
        RECT 24.515 206.195 24.865 206.765 ;
        RECT 25.035 206.025 25.205 206.935 ;
        RECT 25.380 206.670 25.835 207.435 ;
        RECT 26.110 207.055 27.410 207.265 ;
        RECT 27.665 207.075 27.995 207.435 ;
        RECT 27.240 206.905 27.410 207.055 ;
        RECT 28.165 206.935 28.425 207.265 ;
        RECT 26.310 206.445 26.530 206.845 ;
        RECT 25.375 206.245 25.865 206.445 ;
        RECT 26.055 206.235 26.530 206.445 ;
        RECT 26.775 206.445 26.985 206.845 ;
        RECT 27.240 206.780 27.995 206.905 ;
        RECT 27.240 206.735 28.085 206.780 ;
        RECT 27.815 206.615 28.085 206.735 ;
        RECT 26.775 206.235 27.105 206.445 ;
        RECT 27.275 206.175 27.685 206.480 ;
        RECT 24.175 205.855 25.205 206.025 ;
        RECT 23.125 205.515 24.245 205.685 ;
        RECT 23.125 205.055 23.385 205.515 ;
        RECT 23.560 204.885 23.815 205.345 ;
        RECT 23.985 205.055 24.245 205.515 ;
        RECT 24.415 204.885 24.725 205.685 ;
        RECT 24.895 205.055 25.205 205.855 ;
        RECT 25.380 206.005 26.555 206.065 ;
        RECT 27.915 206.040 28.085 206.615 ;
        RECT 27.885 206.005 28.085 206.040 ;
        RECT 25.380 205.895 28.085 206.005 ;
        RECT 25.380 205.275 25.635 205.895 ;
        RECT 26.225 205.835 28.025 205.895 ;
        RECT 26.225 205.805 26.555 205.835 ;
        RECT 28.255 205.735 28.425 206.935 ;
        RECT 25.885 205.635 26.070 205.725 ;
        RECT 26.660 205.635 27.495 205.645 ;
        RECT 25.885 205.435 27.495 205.635 ;
        RECT 25.885 205.395 26.115 205.435 ;
        RECT 25.380 205.055 25.715 205.275 ;
        RECT 26.720 204.885 27.075 205.265 ;
        RECT 27.245 205.055 27.495 205.435 ;
        RECT 27.745 204.885 27.995 205.665 ;
        RECT 28.165 205.055 28.425 205.735 ;
        RECT 28.595 206.975 29.155 207.265 ;
        RECT 29.325 206.975 29.575 207.435 ;
        RECT 28.595 205.605 28.845 206.975 ;
        RECT 30.195 206.805 30.525 207.165 ;
        RECT 29.135 206.615 30.525 206.805 ;
        RECT 30.895 206.665 33.485 207.435 ;
        RECT 34.115 206.710 34.405 207.435 ;
        RECT 34.575 206.935 34.875 207.265 ;
        RECT 35.045 206.955 35.320 207.435 ;
        RECT 29.135 206.525 29.305 206.615 ;
        RECT 29.015 206.195 29.305 206.525 ;
        RECT 29.475 206.195 29.815 206.445 ;
        RECT 30.035 206.195 30.710 206.445 ;
        RECT 29.135 205.945 29.305 206.195 ;
        RECT 29.135 205.775 30.075 205.945 ;
        RECT 30.445 205.835 30.710 206.195 ;
        RECT 30.895 206.145 32.105 206.665 ;
        RECT 32.275 205.975 33.485 206.495 ;
        RECT 28.595 205.055 29.055 205.605 ;
        RECT 29.245 204.885 29.575 205.605 ;
        RECT 29.775 205.225 30.075 205.775 ;
        RECT 30.245 204.885 30.525 205.555 ;
        RECT 30.895 204.885 33.485 205.975 ;
        RECT 34.115 204.885 34.405 206.050 ;
        RECT 34.575 206.025 34.745 206.935 ;
        RECT 35.500 206.785 35.795 207.175 ;
        RECT 35.965 206.955 36.220 207.435 ;
        RECT 36.395 206.785 36.655 207.175 ;
        RECT 36.825 206.955 37.105 207.435 ;
        RECT 37.425 206.885 37.595 207.265 ;
        RECT 37.810 207.055 38.140 207.435 ;
        RECT 34.915 206.195 35.265 206.765 ;
        RECT 35.500 206.615 37.150 206.785 ;
        RECT 37.425 206.715 38.140 206.885 ;
        RECT 35.435 206.275 36.575 206.445 ;
        RECT 35.435 206.025 35.605 206.275 ;
        RECT 36.745 206.105 37.150 206.615 ;
        RECT 37.335 206.165 37.690 206.535 ;
        RECT 37.970 206.525 38.140 206.715 ;
        RECT 38.310 206.690 38.565 207.265 ;
        RECT 37.970 206.195 38.225 206.525 ;
        RECT 34.575 205.855 35.605 206.025 ;
        RECT 36.395 205.935 37.150 206.105 ;
        RECT 37.970 205.985 38.140 206.195 ;
        RECT 34.575 205.055 34.885 205.855 ;
        RECT 36.395 205.685 36.655 205.935 ;
        RECT 37.425 205.815 38.140 205.985 ;
        RECT 38.395 205.960 38.565 206.690 ;
        RECT 38.740 206.595 39.000 207.435 ;
        RECT 39.235 206.955 39.515 207.435 ;
        RECT 39.685 206.785 39.945 207.175 ;
        RECT 40.120 206.955 40.375 207.435 ;
        RECT 40.545 206.785 40.840 207.175 ;
        RECT 41.020 206.955 41.295 207.435 ;
        RECT 41.465 206.935 41.765 207.265 ;
        RECT 39.190 206.615 40.840 206.785 ;
        RECT 39.190 206.105 39.595 206.615 ;
        RECT 39.765 206.275 40.905 206.445 ;
        RECT 35.055 204.885 35.365 205.685 ;
        RECT 35.535 205.515 36.655 205.685 ;
        RECT 35.535 205.055 35.795 205.515 ;
        RECT 35.965 204.885 36.220 205.345 ;
        RECT 36.395 205.055 36.655 205.515 ;
        RECT 36.825 204.885 37.110 205.755 ;
        RECT 37.425 205.055 37.595 205.815 ;
        RECT 37.810 204.885 38.140 205.645 ;
        RECT 38.310 205.055 38.565 205.960 ;
        RECT 38.740 204.885 39.000 206.035 ;
        RECT 39.190 205.935 39.945 206.105 ;
        RECT 39.230 204.885 39.515 205.755 ;
        RECT 39.685 205.685 39.945 205.935 ;
        RECT 40.735 206.025 40.905 206.275 ;
        RECT 41.075 206.195 41.425 206.765 ;
        RECT 41.595 206.025 41.765 206.935 ;
        RECT 41.935 206.685 43.145 207.435 ;
        RECT 40.735 205.855 41.765 206.025 ;
        RECT 39.685 205.515 40.805 205.685 ;
        RECT 39.685 205.055 39.945 205.515 ;
        RECT 40.120 204.885 40.375 205.345 ;
        RECT 40.545 205.055 40.805 205.515 ;
        RECT 40.975 204.885 41.285 205.685 ;
        RECT 41.455 205.055 41.765 205.855 ;
        RECT 41.935 205.975 42.455 206.515 ;
        RECT 42.625 206.145 43.145 206.685 ;
        RECT 41.935 204.885 43.145 205.975 ;
        RECT 8.270 204.715 43.230 204.885 ;
        RECT 8.355 203.625 9.565 204.715 ;
        RECT 9.790 203.845 10.075 204.715 ;
        RECT 10.245 204.085 10.505 204.545 ;
        RECT 10.680 204.255 10.935 204.715 ;
        RECT 11.105 204.085 11.365 204.545 ;
        RECT 10.245 203.915 11.365 204.085 ;
        RECT 11.535 203.915 11.845 204.715 ;
        RECT 10.245 203.665 10.505 203.915 ;
        RECT 12.015 203.745 12.325 204.545 ;
        RECT 8.355 202.915 8.875 203.455 ;
        RECT 9.045 203.085 9.565 203.625 ;
        RECT 9.750 203.495 10.505 203.665 ;
        RECT 11.295 203.575 12.325 203.745 ;
        RECT 9.750 202.985 10.155 203.495 ;
        RECT 11.295 203.325 11.465 203.575 ;
        RECT 10.325 203.155 11.465 203.325 ;
        RECT 8.355 202.165 9.565 202.915 ;
        RECT 9.750 202.815 11.400 202.985 ;
        RECT 11.635 202.835 11.985 203.405 ;
        RECT 9.795 202.165 10.075 202.645 ;
        RECT 10.245 202.425 10.505 202.815 ;
        RECT 10.680 202.165 10.935 202.645 ;
        RECT 11.105 202.425 11.400 202.815 ;
        RECT 12.155 202.665 12.325 203.575 ;
        RECT 11.580 202.165 11.855 202.645 ;
        RECT 12.025 202.335 12.325 202.665 ;
        RECT 12.495 203.640 12.765 204.545 ;
        RECT 12.935 203.955 13.265 204.715 ;
        RECT 13.445 203.785 13.615 204.545 ;
        RECT 12.495 202.840 12.665 203.640 ;
        RECT 12.950 203.615 13.615 203.785 ;
        RECT 13.875 203.865 14.135 204.545 ;
        RECT 14.305 203.935 14.555 204.715 ;
        RECT 14.805 204.165 15.055 204.545 ;
        RECT 15.225 204.335 15.580 204.715 ;
        RECT 16.585 204.325 16.920 204.545 ;
        RECT 16.185 204.165 16.415 204.205 ;
        RECT 14.805 203.965 16.415 204.165 ;
        RECT 14.805 203.955 15.640 203.965 ;
        RECT 16.230 203.875 16.415 203.965 ;
        RECT 12.950 203.470 13.120 203.615 ;
        RECT 12.835 203.140 13.120 203.470 ;
        RECT 12.950 202.885 13.120 203.140 ;
        RECT 13.355 203.065 13.685 203.435 ;
        RECT 12.495 202.335 12.755 202.840 ;
        RECT 12.950 202.715 13.615 202.885 ;
        RECT 12.935 202.165 13.265 202.545 ;
        RECT 13.445 202.335 13.615 202.715 ;
        RECT 13.875 202.675 14.045 203.865 ;
        RECT 15.745 203.765 16.075 203.795 ;
        RECT 14.275 203.705 16.075 203.765 ;
        RECT 16.665 203.705 16.920 204.325 ;
        RECT 17.150 203.845 17.435 204.715 ;
        RECT 17.605 204.085 17.865 204.545 ;
        RECT 18.040 204.255 18.295 204.715 ;
        RECT 18.465 204.085 18.725 204.545 ;
        RECT 17.605 203.915 18.725 204.085 ;
        RECT 18.895 203.915 19.205 204.715 ;
        RECT 14.215 203.595 16.920 203.705 ;
        RECT 17.605 203.665 17.865 203.915 ;
        RECT 18.075 203.865 18.245 203.915 ;
        RECT 19.375 203.745 19.685 204.545 ;
        RECT 14.215 203.560 14.415 203.595 ;
        RECT 14.215 202.985 14.385 203.560 ;
        RECT 15.745 203.535 16.920 203.595 ;
        RECT 17.110 203.495 17.865 203.665 ;
        RECT 18.655 203.575 19.685 203.745 ;
        RECT 19.855 203.625 21.065 204.715 ;
        RECT 14.615 203.120 15.025 203.425 ;
        RECT 15.195 203.155 15.525 203.365 ;
        RECT 14.215 202.865 14.485 202.985 ;
        RECT 14.215 202.820 15.060 202.865 ;
        RECT 14.305 202.695 15.060 202.820 ;
        RECT 15.315 202.755 15.525 203.155 ;
        RECT 15.770 203.155 16.245 203.365 ;
        RECT 16.435 203.155 16.925 203.355 ;
        RECT 15.770 202.755 15.990 203.155 ;
        RECT 17.110 202.985 17.515 203.495 ;
        RECT 18.655 203.325 18.825 203.575 ;
        RECT 17.685 203.155 18.825 203.325 ;
        RECT 13.875 202.665 14.105 202.675 ;
        RECT 13.875 202.335 14.135 202.665 ;
        RECT 14.890 202.545 15.060 202.695 ;
        RECT 14.305 202.165 14.635 202.525 ;
        RECT 14.890 202.335 16.190 202.545 ;
        RECT 16.465 202.165 16.920 202.930 ;
        RECT 17.110 202.815 18.760 202.985 ;
        RECT 18.995 202.835 19.345 203.405 ;
        RECT 17.155 202.165 17.435 202.645 ;
        RECT 17.605 202.425 17.865 202.815 ;
        RECT 18.040 202.165 18.295 202.645 ;
        RECT 18.465 202.425 18.760 202.815 ;
        RECT 19.515 202.665 19.685 203.575 ;
        RECT 18.940 202.165 19.215 202.645 ;
        RECT 19.385 202.335 19.685 202.665 ;
        RECT 19.855 202.915 20.375 203.455 ;
        RECT 20.545 203.085 21.065 203.625 ;
        RECT 21.235 203.550 21.525 204.715 ;
        RECT 21.695 203.575 22.080 204.545 ;
        RECT 22.250 204.255 22.575 204.715 ;
        RECT 23.095 204.085 23.375 204.545 ;
        RECT 22.250 203.865 23.375 204.085 ;
        RECT 19.855 202.165 21.065 202.915 ;
        RECT 21.695 202.905 21.975 203.575 ;
        RECT 22.250 203.405 22.700 203.865 ;
        RECT 23.565 203.695 23.965 204.545 ;
        RECT 24.365 204.255 24.635 204.715 ;
        RECT 24.805 204.085 25.090 204.545 ;
        RECT 22.145 203.075 22.700 203.405 ;
        RECT 22.870 203.135 23.965 203.695 ;
        RECT 22.250 202.965 22.700 203.075 ;
        RECT 21.235 202.165 21.525 202.890 ;
        RECT 21.695 202.335 22.080 202.905 ;
        RECT 22.250 202.795 23.375 202.965 ;
        RECT 22.250 202.165 22.575 202.625 ;
        RECT 23.095 202.335 23.375 202.795 ;
        RECT 23.565 202.335 23.965 203.135 ;
        RECT 24.135 203.865 25.090 204.085 ;
        RECT 24.135 202.965 24.345 203.865 ;
        RECT 24.515 203.135 25.205 203.695 ;
        RECT 25.375 203.625 27.045 204.715 ;
        RECT 24.135 202.795 25.090 202.965 ;
        RECT 24.365 202.165 24.635 202.625 ;
        RECT 24.805 202.335 25.090 202.795 ;
        RECT 25.375 202.935 26.125 203.455 ;
        RECT 26.295 203.105 27.045 203.625 ;
        RECT 27.265 203.575 27.515 204.715 ;
        RECT 27.685 203.525 27.935 204.405 ;
        RECT 28.105 203.575 28.410 204.715 ;
        RECT 28.750 204.335 29.080 204.715 ;
        RECT 29.260 204.165 29.430 204.455 ;
        RECT 29.600 204.255 29.850 204.715 ;
        RECT 28.630 203.995 29.430 204.165 ;
        RECT 30.020 204.205 30.890 204.545 ;
        RECT 25.375 202.165 27.045 202.935 ;
        RECT 27.265 202.165 27.515 202.920 ;
        RECT 27.685 202.875 27.890 203.525 ;
        RECT 28.630 203.405 28.800 203.995 ;
        RECT 30.020 203.825 30.190 204.205 ;
        RECT 31.125 204.085 31.295 204.545 ;
        RECT 31.465 204.255 31.835 204.715 ;
        RECT 32.130 204.115 32.300 204.455 ;
        RECT 32.470 204.285 32.800 204.715 ;
        RECT 33.035 204.115 33.205 204.455 ;
        RECT 28.970 203.655 30.190 203.825 ;
        RECT 30.360 203.745 30.820 204.035 ;
        RECT 31.125 203.915 31.685 204.085 ;
        RECT 32.130 203.945 33.205 204.115 ;
        RECT 33.375 204.215 34.055 204.545 ;
        RECT 34.270 204.215 34.520 204.545 ;
        RECT 34.690 204.255 34.940 204.715 ;
        RECT 31.515 203.775 31.685 203.915 ;
        RECT 30.360 203.735 31.325 203.745 ;
        RECT 30.020 203.565 30.190 203.655 ;
        RECT 30.650 203.575 31.325 203.735 ;
        RECT 28.060 203.375 28.800 203.405 ;
        RECT 28.060 203.075 28.975 203.375 ;
        RECT 28.650 202.900 28.975 203.075 ;
        RECT 27.685 202.345 27.935 202.875 ;
        RECT 28.105 202.165 28.410 202.625 ;
        RECT 28.655 202.545 28.975 202.900 ;
        RECT 29.145 203.115 29.685 203.485 ;
        RECT 30.020 203.395 30.425 203.565 ;
        RECT 29.145 202.715 29.385 203.115 ;
        RECT 29.865 202.945 30.085 203.225 ;
        RECT 29.555 202.775 30.085 202.945 ;
        RECT 29.555 202.545 29.725 202.775 ;
        RECT 30.255 202.615 30.425 203.395 ;
        RECT 30.595 202.785 30.945 203.405 ;
        RECT 31.115 202.785 31.325 203.575 ;
        RECT 31.515 203.605 33.015 203.775 ;
        RECT 31.515 202.915 31.685 203.605 ;
        RECT 33.375 203.435 33.545 204.215 ;
        RECT 34.350 204.085 34.520 204.215 ;
        RECT 31.855 203.265 33.545 203.435 ;
        RECT 33.715 203.655 34.180 204.045 ;
        RECT 34.350 203.915 34.745 204.085 ;
        RECT 31.855 203.085 32.025 203.265 ;
        RECT 28.655 202.375 29.725 202.545 ;
        RECT 29.895 202.165 30.085 202.605 ;
        RECT 30.255 202.335 31.205 202.615 ;
        RECT 31.515 202.525 31.775 202.915 ;
        RECT 32.195 202.845 32.985 203.095 ;
        RECT 31.425 202.355 31.775 202.525 ;
        RECT 31.985 202.165 32.315 202.625 ;
        RECT 33.190 202.555 33.360 203.265 ;
        RECT 33.715 203.065 33.885 203.655 ;
        RECT 33.530 202.845 33.885 203.065 ;
        RECT 34.055 202.845 34.405 203.465 ;
        RECT 34.575 202.555 34.745 203.915 ;
        RECT 35.110 203.745 35.435 204.530 ;
        RECT 34.915 202.695 35.375 203.745 ;
        RECT 33.190 202.385 34.045 202.555 ;
        RECT 34.250 202.385 34.745 202.555 ;
        RECT 34.915 202.165 35.245 202.525 ;
        RECT 35.605 202.425 35.775 204.545 ;
        RECT 35.945 204.215 36.275 204.715 ;
        RECT 36.445 204.045 36.700 204.545 ;
        RECT 35.950 203.875 36.700 204.045 ;
        RECT 35.950 202.885 36.180 203.875 ;
        RECT 36.875 203.865 37.135 204.545 ;
        RECT 37.305 203.935 37.555 204.715 ;
        RECT 37.805 204.165 38.055 204.545 ;
        RECT 38.225 204.335 38.580 204.715 ;
        RECT 39.585 204.325 39.920 204.545 ;
        RECT 39.185 204.165 39.415 204.205 ;
        RECT 37.805 203.965 39.415 204.165 ;
        RECT 37.805 203.955 38.640 203.965 ;
        RECT 39.230 203.875 39.415 203.965 ;
        RECT 36.350 203.055 36.700 203.705 ;
        RECT 35.950 202.715 36.700 202.885 ;
        RECT 35.945 202.165 36.275 202.545 ;
        RECT 36.445 202.425 36.700 202.715 ;
        RECT 36.875 202.665 37.045 203.865 ;
        RECT 38.745 203.765 39.075 203.795 ;
        RECT 37.275 203.705 39.075 203.765 ;
        RECT 39.665 203.705 39.920 204.325 ;
        RECT 37.215 203.595 39.920 203.705 ;
        RECT 40.185 203.785 40.355 204.545 ;
        RECT 40.570 203.955 40.900 204.715 ;
        RECT 40.185 203.615 40.900 203.785 ;
        RECT 41.070 203.640 41.325 204.545 ;
        RECT 37.215 203.560 37.415 203.595 ;
        RECT 37.215 202.985 37.385 203.560 ;
        RECT 38.745 203.535 39.920 203.595 ;
        RECT 37.615 203.120 38.025 203.425 ;
        RECT 38.195 203.155 38.525 203.365 ;
        RECT 37.215 202.865 37.485 202.985 ;
        RECT 37.215 202.820 38.060 202.865 ;
        RECT 37.305 202.695 38.060 202.820 ;
        RECT 38.315 202.755 38.525 203.155 ;
        RECT 38.770 203.155 39.245 203.365 ;
        RECT 39.435 203.155 39.925 203.355 ;
        RECT 38.770 202.755 38.990 203.155 ;
        RECT 40.095 203.065 40.450 203.435 ;
        RECT 40.730 203.405 40.900 203.615 ;
        RECT 40.730 203.075 40.985 203.405 ;
        RECT 36.875 202.335 37.135 202.665 ;
        RECT 37.890 202.545 38.060 202.695 ;
        RECT 37.305 202.165 37.635 202.525 ;
        RECT 37.890 202.335 39.190 202.545 ;
        RECT 39.465 202.165 39.920 202.930 ;
        RECT 40.730 202.885 40.900 203.075 ;
        RECT 41.155 202.910 41.325 203.640 ;
        RECT 41.500 203.565 41.760 204.715 ;
        RECT 41.935 203.625 43.145 204.715 ;
        RECT 41.935 203.085 42.455 203.625 ;
        RECT 40.185 202.715 40.900 202.885 ;
        RECT 40.185 202.335 40.355 202.715 ;
        RECT 40.570 202.165 40.900 202.545 ;
        RECT 41.070 202.335 41.325 202.910 ;
        RECT 41.500 202.165 41.760 203.005 ;
        RECT 42.625 202.915 43.145 203.455 ;
        RECT 41.935 202.165 43.145 202.915 ;
        RECT 8.270 201.995 43.230 202.165 ;
        RECT 8.355 201.245 9.565 201.995 ;
        RECT 9.825 201.445 9.995 201.825 ;
        RECT 10.175 201.615 10.505 201.995 ;
        RECT 9.825 201.275 10.490 201.445 ;
        RECT 10.685 201.320 10.945 201.825 ;
        RECT 8.355 200.705 8.875 201.245 ;
        RECT 9.045 200.535 9.565 201.075 ;
        RECT 9.755 200.725 10.085 201.095 ;
        RECT 10.320 201.020 10.490 201.275 ;
        RECT 10.320 200.690 10.605 201.020 ;
        RECT 10.320 200.545 10.490 200.690 ;
        RECT 8.355 199.445 9.565 200.535 ;
        RECT 9.825 200.375 10.490 200.545 ;
        RECT 10.775 200.520 10.945 201.320 ;
        RECT 9.825 199.615 9.995 200.375 ;
        RECT 10.175 199.445 10.505 200.205 ;
        RECT 10.675 199.615 10.945 200.520 ;
        RECT 11.125 199.625 11.385 201.815 ;
        RECT 11.645 201.625 12.315 201.995 ;
        RECT 12.495 201.445 12.805 201.815 ;
        RECT 11.575 201.245 12.805 201.445 ;
        RECT 11.575 200.575 11.865 201.245 ;
        RECT 12.985 201.065 13.215 201.705 ;
        RECT 13.395 201.265 13.685 201.995 ;
        RECT 13.925 201.240 14.175 201.995 ;
        RECT 14.345 201.285 14.595 201.815 ;
        RECT 14.765 201.535 15.070 201.995 ;
        RECT 15.315 201.615 16.385 201.785 ;
        RECT 12.045 200.755 12.510 201.065 ;
        RECT 12.690 200.755 13.215 201.065 ;
        RECT 13.395 200.755 13.695 201.085 ;
        RECT 14.345 200.635 14.550 201.285 ;
        RECT 15.315 201.260 15.635 201.615 ;
        RECT 15.310 201.085 15.635 201.260 ;
        RECT 14.720 200.785 15.635 201.085 ;
        RECT 15.805 201.045 16.045 201.445 ;
        RECT 16.215 201.385 16.385 201.615 ;
        RECT 16.555 201.555 16.745 201.995 ;
        RECT 16.915 201.545 17.865 201.825 ;
        RECT 18.085 201.635 18.435 201.805 ;
        RECT 16.215 201.215 16.745 201.385 ;
        RECT 14.720 200.755 15.460 200.785 ;
        RECT 11.575 200.355 12.345 200.575 ;
        RECT 11.555 199.445 11.895 200.175 ;
        RECT 12.075 199.625 12.345 200.355 ;
        RECT 12.525 200.335 13.685 200.575 ;
        RECT 12.525 199.625 12.755 200.335 ;
        RECT 12.925 199.445 13.255 200.155 ;
        RECT 13.425 199.625 13.685 200.335 ;
        RECT 13.925 199.445 14.175 200.585 ;
        RECT 14.345 199.755 14.595 200.635 ;
        RECT 14.765 199.445 15.070 200.585 ;
        RECT 15.290 200.165 15.460 200.755 ;
        RECT 15.805 200.675 16.345 201.045 ;
        RECT 16.525 200.935 16.745 201.215 ;
        RECT 16.915 200.765 17.085 201.545 ;
        RECT 16.680 200.595 17.085 200.765 ;
        RECT 17.255 200.755 17.605 201.375 ;
        RECT 16.680 200.505 16.850 200.595 ;
        RECT 17.775 200.585 17.985 201.375 ;
        RECT 15.630 200.335 16.850 200.505 ;
        RECT 17.310 200.425 17.985 200.585 ;
        RECT 15.290 199.995 16.090 200.165 ;
        RECT 15.410 199.445 15.740 199.825 ;
        RECT 15.920 199.705 16.090 199.995 ;
        RECT 16.680 199.955 16.850 200.335 ;
        RECT 17.020 200.415 17.985 200.425 ;
        RECT 18.175 201.245 18.435 201.635 ;
        RECT 18.645 201.535 18.975 201.995 ;
        RECT 19.850 201.605 20.705 201.775 ;
        RECT 20.910 201.605 21.405 201.775 ;
        RECT 21.575 201.635 21.905 201.995 ;
        RECT 18.175 200.555 18.345 201.245 ;
        RECT 18.515 200.895 18.685 201.075 ;
        RECT 18.855 201.065 19.645 201.315 ;
        RECT 19.850 200.895 20.020 201.605 ;
        RECT 20.190 201.095 20.545 201.315 ;
        RECT 18.515 200.725 20.205 200.895 ;
        RECT 17.020 200.125 17.480 200.415 ;
        RECT 18.175 200.385 19.675 200.555 ;
        RECT 18.175 200.245 18.345 200.385 ;
        RECT 17.785 200.075 18.345 200.245 ;
        RECT 16.260 199.445 16.510 199.905 ;
        RECT 16.680 199.615 17.550 199.955 ;
        RECT 17.785 199.615 17.955 200.075 ;
        RECT 18.790 200.045 19.865 200.215 ;
        RECT 18.125 199.445 18.495 199.905 ;
        RECT 18.790 199.705 18.960 200.045 ;
        RECT 19.130 199.445 19.460 199.875 ;
        RECT 19.695 199.705 19.865 200.045 ;
        RECT 20.035 199.945 20.205 200.725 ;
        RECT 20.375 200.505 20.545 201.095 ;
        RECT 20.715 200.695 21.065 201.315 ;
        RECT 20.375 200.115 20.840 200.505 ;
        RECT 21.235 200.245 21.405 201.605 ;
        RECT 21.575 200.415 22.035 201.465 ;
        RECT 21.010 200.075 21.405 200.245 ;
        RECT 21.010 199.945 21.180 200.075 ;
        RECT 20.035 199.615 20.715 199.945 ;
        RECT 20.930 199.615 21.180 199.945 ;
        RECT 21.350 199.445 21.600 199.905 ;
        RECT 21.770 199.630 22.095 200.415 ;
        RECT 22.265 199.615 22.435 201.735 ;
        RECT 22.605 201.615 22.935 201.995 ;
        RECT 23.105 201.445 23.360 201.735 ;
        RECT 22.610 201.275 23.360 201.445 ;
        RECT 22.610 200.285 22.840 201.275 ;
        RECT 23.535 201.245 24.745 201.995 ;
        RECT 25.005 201.445 25.175 201.825 ;
        RECT 25.355 201.615 25.685 201.995 ;
        RECT 25.005 201.275 25.670 201.445 ;
        RECT 25.865 201.320 26.125 201.825 ;
        RECT 23.010 200.455 23.360 201.105 ;
        RECT 23.535 200.705 24.055 201.245 ;
        RECT 24.225 200.535 24.745 201.075 ;
        RECT 24.935 200.725 25.265 201.095 ;
        RECT 25.500 201.020 25.670 201.275 ;
        RECT 25.500 200.690 25.785 201.020 ;
        RECT 25.500 200.545 25.670 200.690 ;
        RECT 22.610 200.115 23.360 200.285 ;
        RECT 22.605 199.445 22.935 199.945 ;
        RECT 23.105 199.615 23.360 200.115 ;
        RECT 23.535 199.445 24.745 200.535 ;
        RECT 25.005 200.375 25.670 200.545 ;
        RECT 25.955 200.520 26.125 201.320 ;
        RECT 25.005 199.615 25.175 200.375 ;
        RECT 25.355 199.445 25.685 200.205 ;
        RECT 25.855 199.615 26.125 200.520 ;
        RECT 26.295 201.255 26.680 201.825 ;
        RECT 26.850 201.535 27.175 201.995 ;
        RECT 27.695 201.365 27.975 201.825 ;
        RECT 26.295 200.585 26.575 201.255 ;
        RECT 26.850 201.195 27.975 201.365 ;
        RECT 26.850 201.085 27.300 201.195 ;
        RECT 26.745 200.755 27.300 201.085 ;
        RECT 28.165 201.025 28.565 201.825 ;
        RECT 28.965 201.535 29.235 201.995 ;
        RECT 29.405 201.365 29.690 201.825 ;
        RECT 26.295 199.615 26.680 200.585 ;
        RECT 26.850 200.295 27.300 200.755 ;
        RECT 27.470 200.465 28.565 201.025 ;
        RECT 26.850 200.075 27.975 200.295 ;
        RECT 26.850 199.445 27.175 199.905 ;
        RECT 27.695 199.615 27.975 200.075 ;
        RECT 28.165 199.615 28.565 200.465 ;
        RECT 28.735 201.195 29.690 201.365 ;
        RECT 30.090 201.365 30.375 201.825 ;
        RECT 30.545 201.535 30.815 201.995 ;
        RECT 30.090 201.195 31.045 201.365 ;
        RECT 28.735 200.295 28.945 201.195 ;
        RECT 29.115 200.465 29.805 201.025 ;
        RECT 29.975 200.465 30.665 201.025 ;
        RECT 30.835 200.295 31.045 201.195 ;
        RECT 28.735 200.075 29.690 200.295 ;
        RECT 28.965 199.445 29.235 199.905 ;
        RECT 29.405 199.615 29.690 200.075 ;
        RECT 30.090 200.075 31.045 200.295 ;
        RECT 31.215 201.025 31.615 201.825 ;
        RECT 31.805 201.365 32.085 201.825 ;
        RECT 32.605 201.535 32.930 201.995 ;
        RECT 31.805 201.195 32.930 201.365 ;
        RECT 33.100 201.255 33.485 201.825 ;
        RECT 34.115 201.270 34.405 201.995 ;
        RECT 32.480 201.085 32.930 201.195 ;
        RECT 31.215 200.465 32.310 201.025 ;
        RECT 32.480 200.755 33.035 201.085 ;
        RECT 30.090 199.615 30.375 200.075 ;
        RECT 30.545 199.445 30.815 199.905 ;
        RECT 31.215 199.615 31.615 200.465 ;
        RECT 32.480 200.295 32.930 200.755 ;
        RECT 33.205 200.585 33.485 201.255 ;
        RECT 34.575 201.255 34.960 201.825 ;
        RECT 35.130 201.535 35.455 201.995 ;
        RECT 35.975 201.365 36.255 201.825 ;
        RECT 31.805 200.075 32.930 200.295 ;
        RECT 31.805 199.615 32.085 200.075 ;
        RECT 32.605 199.445 32.930 199.905 ;
        RECT 33.100 199.615 33.485 200.585 ;
        RECT 34.115 199.445 34.405 200.610 ;
        RECT 34.575 200.585 34.855 201.255 ;
        RECT 35.130 201.195 36.255 201.365 ;
        RECT 35.130 201.085 35.580 201.195 ;
        RECT 35.025 200.755 35.580 201.085 ;
        RECT 36.445 201.025 36.845 201.825 ;
        RECT 37.245 201.535 37.515 201.995 ;
        RECT 37.685 201.365 37.970 201.825 ;
        RECT 34.575 199.615 34.960 200.585 ;
        RECT 35.130 200.295 35.580 200.755 ;
        RECT 35.750 200.465 36.845 201.025 ;
        RECT 35.130 200.075 36.255 200.295 ;
        RECT 35.130 199.445 35.455 199.905 ;
        RECT 35.975 199.615 36.255 200.075 ;
        RECT 36.445 199.615 36.845 200.465 ;
        RECT 37.015 201.195 37.970 201.365 ;
        RECT 38.255 201.495 38.515 201.825 ;
        RECT 38.685 201.635 39.015 201.995 ;
        RECT 39.270 201.615 40.570 201.825 ;
        RECT 38.255 201.485 38.485 201.495 ;
        RECT 37.015 200.295 37.225 201.195 ;
        RECT 37.395 200.465 38.085 201.025 ;
        RECT 38.255 200.295 38.425 201.485 ;
        RECT 39.270 201.465 39.440 201.615 ;
        RECT 38.685 201.340 39.440 201.465 ;
        RECT 38.595 201.295 39.440 201.340 ;
        RECT 38.595 201.175 38.865 201.295 ;
        RECT 38.595 200.600 38.765 201.175 ;
        RECT 38.995 200.735 39.405 201.040 ;
        RECT 39.695 201.005 39.905 201.405 ;
        RECT 39.575 200.795 39.905 201.005 ;
        RECT 40.150 201.005 40.370 201.405 ;
        RECT 40.845 201.230 41.300 201.995 ;
        RECT 41.935 201.245 43.145 201.995 ;
        RECT 40.150 200.795 40.625 201.005 ;
        RECT 40.815 200.805 41.305 201.005 ;
        RECT 38.595 200.565 38.795 200.600 ;
        RECT 40.125 200.565 41.300 200.625 ;
        RECT 38.595 200.455 41.300 200.565 ;
        RECT 38.655 200.395 40.455 200.455 ;
        RECT 40.125 200.365 40.455 200.395 ;
        RECT 37.015 200.075 37.970 200.295 ;
        RECT 37.245 199.445 37.515 199.905 ;
        RECT 37.685 199.615 37.970 200.075 ;
        RECT 38.255 199.615 38.515 200.295 ;
        RECT 38.685 199.445 38.935 200.225 ;
        RECT 39.185 200.195 40.020 200.205 ;
        RECT 40.610 200.195 40.795 200.285 ;
        RECT 39.185 199.995 40.795 200.195 ;
        RECT 39.185 199.615 39.435 199.995 ;
        RECT 40.565 199.955 40.795 199.995 ;
        RECT 41.045 199.835 41.300 200.455 ;
        RECT 39.605 199.445 39.960 199.825 ;
        RECT 40.965 199.615 41.300 199.835 ;
        RECT 41.935 200.535 42.455 201.075 ;
        RECT 42.625 200.705 43.145 201.245 ;
        RECT 41.935 199.445 43.145 200.535 ;
        RECT 8.270 199.275 43.230 199.445 ;
        RECT 8.355 198.185 9.565 199.275 ;
        RECT 8.355 197.475 8.875 198.015 ;
        RECT 9.045 197.645 9.565 198.185 ;
        RECT 9.735 198.305 10.045 199.105 ;
        RECT 10.215 198.475 10.525 199.275 ;
        RECT 10.695 198.645 10.955 199.105 ;
        RECT 11.125 198.815 11.380 199.275 ;
        RECT 11.555 198.645 11.815 199.105 ;
        RECT 10.695 198.475 11.815 198.645 ;
        RECT 11.175 198.425 11.345 198.475 ;
        RECT 9.735 198.135 10.765 198.305 ;
        RECT 8.355 196.725 9.565 197.475 ;
        RECT 9.735 197.225 9.905 198.135 ;
        RECT 10.075 197.395 10.425 197.965 ;
        RECT 10.595 197.885 10.765 198.135 ;
        RECT 11.555 198.225 11.815 198.475 ;
        RECT 11.985 198.405 12.270 199.275 ;
        RECT 12.550 198.405 12.835 199.275 ;
        RECT 13.005 198.645 13.265 199.105 ;
        RECT 13.440 198.815 13.695 199.275 ;
        RECT 13.865 198.645 14.125 199.105 ;
        RECT 13.005 198.475 14.125 198.645 ;
        RECT 14.295 198.475 14.605 199.275 ;
        RECT 13.005 198.225 13.265 198.475 ;
        RECT 14.775 198.305 15.085 199.105 ;
        RECT 11.555 198.055 12.310 198.225 ;
        RECT 10.595 197.715 11.735 197.885 ;
        RECT 11.905 197.545 12.310 198.055 ;
        RECT 10.660 197.375 12.310 197.545 ;
        RECT 12.510 198.055 13.265 198.225 ;
        RECT 14.055 198.135 15.085 198.305 ;
        RECT 12.510 197.545 12.915 198.055 ;
        RECT 14.055 197.885 14.225 198.135 ;
        RECT 13.085 197.715 14.225 197.885 ;
        RECT 12.510 197.375 14.160 197.545 ;
        RECT 14.395 197.395 14.745 197.965 ;
        RECT 9.735 196.895 10.035 197.225 ;
        RECT 10.205 196.725 10.480 197.205 ;
        RECT 10.660 196.985 10.955 197.375 ;
        RECT 11.125 196.725 11.380 197.205 ;
        RECT 11.555 196.985 11.815 197.375 ;
        RECT 11.985 196.725 12.265 197.205 ;
        RECT 12.555 196.725 12.835 197.205 ;
        RECT 13.005 196.985 13.265 197.375 ;
        RECT 13.440 196.725 13.695 197.205 ;
        RECT 13.865 196.985 14.160 197.375 ;
        RECT 14.915 197.225 15.085 198.135 ;
        RECT 15.260 198.885 15.595 199.105 ;
        RECT 16.600 198.895 16.955 199.275 ;
        RECT 15.260 198.265 15.515 198.885 ;
        RECT 15.765 198.725 15.995 198.765 ;
        RECT 17.125 198.725 17.375 199.105 ;
        RECT 15.765 198.525 17.375 198.725 ;
        RECT 15.765 198.435 15.950 198.525 ;
        RECT 16.540 198.515 17.375 198.525 ;
        RECT 17.625 198.495 17.875 199.275 ;
        RECT 18.045 198.425 18.305 199.105 ;
        RECT 16.105 198.325 16.435 198.355 ;
        RECT 16.105 198.265 17.905 198.325 ;
        RECT 15.260 198.155 17.965 198.265 ;
        RECT 15.260 198.095 16.435 198.155 ;
        RECT 17.765 198.120 17.965 198.155 ;
        RECT 15.255 197.715 15.745 197.915 ;
        RECT 15.935 197.715 16.410 197.925 ;
        RECT 14.340 196.725 14.615 197.205 ;
        RECT 14.785 196.895 15.085 197.225 ;
        RECT 15.260 196.725 15.715 197.490 ;
        RECT 16.190 197.315 16.410 197.715 ;
        RECT 16.655 197.715 16.985 197.925 ;
        RECT 16.655 197.315 16.865 197.715 ;
        RECT 17.155 197.680 17.565 197.985 ;
        RECT 17.795 197.545 17.965 198.120 ;
        RECT 17.695 197.425 17.965 197.545 ;
        RECT 17.120 197.380 17.965 197.425 ;
        RECT 17.120 197.255 17.875 197.380 ;
        RECT 17.120 197.105 17.290 197.255 ;
        RECT 18.135 197.235 18.305 198.425 ;
        RECT 18.530 198.405 18.815 199.275 ;
        RECT 18.985 198.645 19.245 199.105 ;
        RECT 19.420 198.815 19.675 199.275 ;
        RECT 19.845 198.645 20.105 199.105 ;
        RECT 18.985 198.475 20.105 198.645 ;
        RECT 20.275 198.475 20.585 199.275 ;
        RECT 18.985 198.225 19.245 198.475 ;
        RECT 20.755 198.305 21.065 199.105 ;
        RECT 18.490 198.055 19.245 198.225 ;
        RECT 20.035 198.135 21.065 198.305 ;
        RECT 18.490 197.545 18.895 198.055 ;
        RECT 20.035 197.885 20.205 198.135 ;
        RECT 19.065 197.715 20.205 197.885 ;
        RECT 18.490 197.375 20.140 197.545 ;
        RECT 20.375 197.395 20.725 197.965 ;
        RECT 18.075 197.225 18.305 197.235 ;
        RECT 15.990 196.895 17.290 197.105 ;
        RECT 17.545 196.725 17.875 197.085 ;
        RECT 18.045 196.895 18.305 197.225 ;
        RECT 18.535 196.725 18.815 197.205 ;
        RECT 18.985 196.985 19.245 197.375 ;
        RECT 19.420 196.725 19.675 197.205 ;
        RECT 19.845 196.985 20.140 197.375 ;
        RECT 20.895 197.225 21.065 198.135 ;
        RECT 21.235 198.110 21.525 199.275 ;
        RECT 20.320 196.725 20.595 197.205 ;
        RECT 20.765 196.895 21.065 197.225 ;
        RECT 21.235 196.725 21.525 197.450 ;
        RECT 21.705 196.905 21.965 199.095 ;
        RECT 22.135 198.545 22.475 199.275 ;
        RECT 22.655 198.365 22.925 199.095 ;
        RECT 22.155 198.145 22.925 198.365 ;
        RECT 23.105 198.385 23.335 199.095 ;
        RECT 23.505 198.565 23.835 199.275 ;
        RECT 24.005 198.385 24.265 199.095 ;
        RECT 23.105 198.145 24.265 198.385 ;
        RECT 24.455 198.185 27.965 199.275 ;
        RECT 22.155 197.475 22.445 198.145 ;
        RECT 22.625 197.655 23.090 197.965 ;
        RECT 23.270 197.655 23.795 197.965 ;
        RECT 22.155 197.275 23.385 197.475 ;
        RECT 22.225 196.725 22.895 197.095 ;
        RECT 23.075 196.905 23.385 197.275 ;
        RECT 23.565 197.015 23.795 197.655 ;
        RECT 23.975 197.635 24.275 197.965 ;
        RECT 24.455 197.495 26.105 198.015 ;
        RECT 26.275 197.665 27.965 198.185 ;
        RECT 29.055 198.200 29.325 199.105 ;
        RECT 29.495 198.515 29.825 199.275 ;
        RECT 30.005 198.345 30.175 199.105 ;
        RECT 23.975 196.725 24.265 197.455 ;
        RECT 24.455 196.725 27.965 197.495 ;
        RECT 29.055 197.400 29.225 198.200 ;
        RECT 29.510 198.175 30.175 198.345 ;
        RECT 29.510 198.030 29.680 198.175 ;
        RECT 30.485 198.135 30.735 199.275 ;
        RECT 29.395 197.700 29.680 198.030 ;
        RECT 30.905 198.085 31.155 198.965 ;
        RECT 31.325 198.135 31.630 199.275 ;
        RECT 31.970 198.895 32.300 199.275 ;
        RECT 32.480 198.725 32.650 199.015 ;
        RECT 32.820 198.815 33.070 199.275 ;
        RECT 31.850 198.555 32.650 198.725 ;
        RECT 33.240 198.765 34.110 199.105 ;
        RECT 29.510 197.445 29.680 197.700 ;
        RECT 29.915 197.625 30.245 197.995 ;
        RECT 29.055 196.895 29.315 197.400 ;
        RECT 29.510 197.275 30.175 197.445 ;
        RECT 29.495 196.725 29.825 197.105 ;
        RECT 30.005 196.895 30.175 197.275 ;
        RECT 30.485 196.725 30.735 197.480 ;
        RECT 30.905 197.435 31.110 198.085 ;
        RECT 31.850 197.965 32.020 198.555 ;
        RECT 33.240 198.385 33.410 198.765 ;
        RECT 34.345 198.645 34.515 199.105 ;
        RECT 34.685 198.815 35.055 199.275 ;
        RECT 35.350 198.675 35.520 199.015 ;
        RECT 35.690 198.845 36.020 199.275 ;
        RECT 36.255 198.675 36.425 199.015 ;
        RECT 32.190 198.215 33.410 198.385 ;
        RECT 33.580 198.305 34.040 198.595 ;
        RECT 34.345 198.475 34.905 198.645 ;
        RECT 35.350 198.505 36.425 198.675 ;
        RECT 36.595 198.775 37.275 199.105 ;
        RECT 37.490 198.775 37.740 199.105 ;
        RECT 37.910 198.815 38.160 199.275 ;
        RECT 34.735 198.335 34.905 198.475 ;
        RECT 33.580 198.295 34.545 198.305 ;
        RECT 33.240 198.125 33.410 198.215 ;
        RECT 33.870 198.135 34.545 198.295 ;
        RECT 31.280 197.935 32.020 197.965 ;
        RECT 31.280 197.635 32.195 197.935 ;
        RECT 31.870 197.460 32.195 197.635 ;
        RECT 30.905 196.905 31.155 197.435 ;
        RECT 31.325 196.725 31.630 197.185 ;
        RECT 31.875 197.105 32.195 197.460 ;
        RECT 32.365 197.675 32.905 198.045 ;
        RECT 33.240 197.955 33.645 198.125 ;
        RECT 32.365 197.275 32.605 197.675 ;
        RECT 33.085 197.505 33.305 197.785 ;
        RECT 32.775 197.335 33.305 197.505 ;
        RECT 32.775 197.105 32.945 197.335 ;
        RECT 33.475 197.175 33.645 197.955 ;
        RECT 33.815 197.345 34.165 197.965 ;
        RECT 34.335 197.345 34.545 198.135 ;
        RECT 34.735 198.165 36.235 198.335 ;
        RECT 34.735 197.475 34.905 198.165 ;
        RECT 36.595 197.995 36.765 198.775 ;
        RECT 37.570 198.645 37.740 198.775 ;
        RECT 35.075 197.825 36.765 197.995 ;
        RECT 36.935 198.215 37.400 198.605 ;
        RECT 37.570 198.475 37.965 198.645 ;
        RECT 35.075 197.645 35.245 197.825 ;
        RECT 31.875 196.935 32.945 197.105 ;
        RECT 33.115 196.725 33.305 197.165 ;
        RECT 33.475 196.895 34.425 197.175 ;
        RECT 34.735 197.085 34.995 197.475 ;
        RECT 35.415 197.405 36.205 197.655 ;
        RECT 34.645 196.915 34.995 197.085 ;
        RECT 35.205 196.725 35.535 197.185 ;
        RECT 36.410 197.115 36.580 197.825 ;
        RECT 36.935 197.625 37.105 198.215 ;
        RECT 36.750 197.405 37.105 197.625 ;
        RECT 37.275 197.405 37.625 198.025 ;
        RECT 37.795 197.115 37.965 198.475 ;
        RECT 38.330 198.305 38.655 199.090 ;
        RECT 38.135 197.255 38.595 198.305 ;
        RECT 36.410 196.945 37.265 197.115 ;
        RECT 37.470 196.945 37.965 197.115 ;
        RECT 38.135 196.725 38.465 197.085 ;
        RECT 38.825 196.985 38.995 199.105 ;
        RECT 39.165 198.775 39.495 199.275 ;
        RECT 39.665 198.605 39.920 199.105 ;
        RECT 39.170 198.435 39.920 198.605 ;
        RECT 39.170 197.445 39.400 198.435 ;
        RECT 39.570 197.615 39.920 198.265 ;
        RECT 40.095 198.185 41.765 199.275 ;
        RECT 40.095 197.495 40.845 198.015 ;
        RECT 41.015 197.665 41.765 198.185 ;
        RECT 41.935 198.185 43.145 199.275 ;
        RECT 41.935 197.645 42.455 198.185 ;
        RECT 39.170 197.275 39.920 197.445 ;
        RECT 39.165 196.725 39.495 197.105 ;
        RECT 39.665 196.985 39.920 197.275 ;
        RECT 40.095 196.725 41.765 197.495 ;
        RECT 42.625 197.475 43.145 198.015 ;
        RECT 41.935 196.725 43.145 197.475 ;
        RECT 8.270 196.555 43.230 196.725 ;
        RECT 8.355 195.805 9.565 196.555 ;
        RECT 9.735 196.095 10.295 196.385 ;
        RECT 10.465 196.095 10.715 196.555 ;
        RECT 8.355 195.265 8.875 195.805 ;
        RECT 9.045 195.095 9.565 195.635 ;
        RECT 8.355 194.005 9.565 195.095 ;
        RECT 9.735 194.725 9.985 196.095 ;
        RECT 11.335 195.925 11.665 196.285 ;
        RECT 10.275 195.735 11.665 195.925 ;
        RECT 12.125 196.005 12.295 196.295 ;
        RECT 12.465 196.175 12.795 196.555 ;
        RECT 12.125 195.835 12.790 196.005 ;
        RECT 10.275 195.645 10.445 195.735 ;
        RECT 10.155 195.315 10.445 195.645 ;
        RECT 10.615 195.315 10.955 195.565 ;
        RECT 11.175 195.315 11.850 195.565 ;
        RECT 10.275 195.065 10.445 195.315 ;
        RECT 10.275 194.895 11.215 195.065 ;
        RECT 11.585 194.955 11.850 195.315 ;
        RECT 12.040 195.015 12.390 195.665 ;
        RECT 9.735 194.175 10.195 194.725 ;
        RECT 10.385 194.005 10.715 194.725 ;
        RECT 10.915 194.345 11.215 194.895 ;
        RECT 12.560 194.845 12.790 195.835 ;
        RECT 12.125 194.675 12.790 194.845 ;
        RECT 11.385 194.005 11.665 194.675 ;
        RECT 12.125 194.175 12.295 194.675 ;
        RECT 12.465 194.005 12.795 194.505 ;
        RECT 12.965 194.175 13.190 196.295 ;
        RECT 13.405 196.175 13.735 196.555 ;
        RECT 13.905 196.005 14.075 196.335 ;
        RECT 14.375 196.175 15.390 196.375 ;
        RECT 13.380 195.815 14.075 196.005 ;
        RECT 13.380 194.845 13.550 195.815 ;
        RECT 13.720 195.015 14.130 195.635 ;
        RECT 14.300 195.065 14.520 195.935 ;
        RECT 14.700 195.625 15.050 195.995 ;
        RECT 15.220 195.445 15.390 196.175 ;
        RECT 15.560 196.115 15.970 196.555 ;
        RECT 16.260 195.915 16.510 196.345 ;
        RECT 16.710 196.095 17.030 196.555 ;
        RECT 17.590 196.165 18.440 196.335 ;
        RECT 15.560 195.575 15.970 195.905 ;
        RECT 16.260 195.575 16.680 195.915 ;
        RECT 14.970 195.405 15.390 195.445 ;
        RECT 14.970 195.235 16.320 195.405 ;
        RECT 13.380 194.675 14.075 194.845 ;
        RECT 14.300 194.685 14.800 195.065 ;
        RECT 13.405 194.005 13.735 194.505 ;
        RECT 13.905 194.175 14.075 194.675 ;
        RECT 14.970 194.390 15.140 195.235 ;
        RECT 16.070 195.075 16.320 195.235 ;
        RECT 15.310 194.805 15.560 195.065 ;
        RECT 16.490 194.805 16.680 195.575 ;
        RECT 15.310 194.555 16.680 194.805 ;
        RECT 16.850 195.745 18.100 195.915 ;
        RECT 16.850 194.985 17.020 195.745 ;
        RECT 17.770 195.625 18.100 195.745 ;
        RECT 17.190 195.165 17.370 195.575 ;
        RECT 18.270 195.405 18.440 196.165 ;
        RECT 18.640 196.075 19.300 196.555 ;
        RECT 19.480 195.960 19.800 196.290 ;
        RECT 18.630 195.635 19.290 195.905 ;
        RECT 18.630 195.575 18.960 195.635 ;
        RECT 19.110 195.405 19.440 195.465 ;
        RECT 17.540 195.235 19.440 195.405 ;
        RECT 16.850 194.675 17.370 194.985 ;
        RECT 17.540 194.725 17.710 195.235 ;
        RECT 19.610 195.065 19.800 195.960 ;
        RECT 17.880 194.895 19.800 195.065 ;
        RECT 19.480 194.875 19.800 194.895 ;
        RECT 20.000 195.645 20.250 196.295 ;
        RECT 20.430 196.095 20.715 196.555 ;
        RECT 20.895 196.215 21.150 196.375 ;
        RECT 20.895 196.045 21.235 196.215 ;
        RECT 20.895 195.845 21.150 196.045 ;
        RECT 20.000 195.315 20.800 195.645 ;
        RECT 17.540 194.555 18.750 194.725 ;
        RECT 14.310 194.220 15.140 194.390 ;
        RECT 15.380 194.005 15.760 194.385 ;
        RECT 15.940 194.265 16.110 194.555 ;
        RECT 17.540 194.475 17.710 194.555 ;
        RECT 16.280 194.005 16.610 194.385 ;
        RECT 17.080 194.225 17.710 194.475 ;
        RECT 17.890 194.005 18.310 194.385 ;
        RECT 18.510 194.265 18.750 194.555 ;
        RECT 18.980 194.005 19.310 194.695 ;
        RECT 19.480 194.265 19.650 194.875 ;
        RECT 20.000 194.725 20.250 195.315 ;
        RECT 20.970 194.985 21.150 195.845 ;
        RECT 21.700 196.005 21.955 196.295 ;
        RECT 22.125 196.175 22.455 196.555 ;
        RECT 21.700 195.835 22.450 196.005 ;
        RECT 21.700 195.015 22.050 195.665 ;
        RECT 19.920 194.215 20.250 194.725 ;
        RECT 20.430 194.005 20.715 194.805 ;
        RECT 20.895 194.315 21.150 194.985 ;
        RECT 22.220 194.845 22.450 195.835 ;
        RECT 21.700 194.675 22.450 194.845 ;
        RECT 21.700 194.175 21.955 194.675 ;
        RECT 22.125 194.005 22.455 194.505 ;
        RECT 22.625 194.175 22.795 196.295 ;
        RECT 23.155 196.195 23.485 196.555 ;
        RECT 23.655 196.165 24.150 196.335 ;
        RECT 24.355 196.165 25.210 196.335 ;
        RECT 23.025 194.975 23.485 196.025 ;
        RECT 22.965 194.190 23.290 194.975 ;
        RECT 23.655 194.805 23.825 196.165 ;
        RECT 23.995 195.255 24.345 195.875 ;
        RECT 24.515 195.655 24.870 195.875 ;
        RECT 24.515 195.065 24.685 195.655 ;
        RECT 25.040 195.455 25.210 196.165 ;
        RECT 26.085 196.095 26.415 196.555 ;
        RECT 26.625 196.195 26.975 196.365 ;
        RECT 25.415 195.625 26.205 195.875 ;
        RECT 26.625 195.805 26.885 196.195 ;
        RECT 27.195 196.105 28.145 196.385 ;
        RECT 28.315 196.115 28.505 196.555 ;
        RECT 28.675 196.175 29.745 196.345 ;
        RECT 26.375 195.455 26.545 195.635 ;
        RECT 23.655 194.635 24.050 194.805 ;
        RECT 24.220 194.675 24.685 195.065 ;
        RECT 24.855 195.285 26.545 195.455 ;
        RECT 23.880 194.505 24.050 194.635 ;
        RECT 24.855 194.505 25.025 195.285 ;
        RECT 26.715 195.115 26.885 195.805 ;
        RECT 25.385 194.945 26.885 195.115 ;
        RECT 27.075 195.145 27.285 195.935 ;
        RECT 27.455 195.315 27.805 195.935 ;
        RECT 27.975 195.325 28.145 196.105 ;
        RECT 28.675 195.945 28.845 196.175 ;
        RECT 28.315 195.775 28.845 195.945 ;
        RECT 28.315 195.495 28.535 195.775 ;
        RECT 29.015 195.605 29.255 196.005 ;
        RECT 27.975 195.155 28.380 195.325 ;
        RECT 28.715 195.235 29.255 195.605 ;
        RECT 29.425 195.820 29.745 196.175 ;
        RECT 29.990 196.095 30.295 196.555 ;
        RECT 30.465 195.845 30.715 196.375 ;
        RECT 29.425 195.645 29.750 195.820 ;
        RECT 29.425 195.345 30.340 195.645 ;
        RECT 29.600 195.315 30.340 195.345 ;
        RECT 27.075 194.985 27.750 195.145 ;
        RECT 28.210 195.065 28.380 195.155 ;
        RECT 27.075 194.975 28.040 194.985 ;
        RECT 26.715 194.805 26.885 194.945 ;
        RECT 23.460 194.005 23.710 194.465 ;
        RECT 23.880 194.175 24.130 194.505 ;
        RECT 24.345 194.175 25.025 194.505 ;
        RECT 25.195 194.605 26.270 194.775 ;
        RECT 26.715 194.635 27.275 194.805 ;
        RECT 27.580 194.685 28.040 194.975 ;
        RECT 28.210 194.895 29.430 195.065 ;
        RECT 25.195 194.265 25.365 194.605 ;
        RECT 25.600 194.005 25.930 194.435 ;
        RECT 26.100 194.265 26.270 194.605 ;
        RECT 26.565 194.005 26.935 194.465 ;
        RECT 27.105 194.175 27.275 194.635 ;
        RECT 28.210 194.515 28.380 194.895 ;
        RECT 29.600 194.725 29.770 195.315 ;
        RECT 30.510 195.195 30.715 195.845 ;
        RECT 30.885 195.800 31.135 196.555 ;
        RECT 31.355 196.055 31.655 196.385 ;
        RECT 31.825 196.075 32.100 196.555 ;
        RECT 27.510 194.175 28.380 194.515 ;
        RECT 28.970 194.555 29.770 194.725 ;
        RECT 28.550 194.005 28.800 194.465 ;
        RECT 28.970 194.265 29.140 194.555 ;
        RECT 29.320 194.005 29.650 194.385 ;
        RECT 29.990 194.005 30.295 195.145 ;
        RECT 30.465 194.315 30.715 195.195 ;
        RECT 31.355 195.145 31.525 196.055 ;
        RECT 32.280 195.905 32.575 196.295 ;
        RECT 32.745 196.075 33.000 196.555 ;
        RECT 33.175 195.905 33.435 196.295 ;
        RECT 33.605 196.075 33.885 196.555 ;
        RECT 31.695 195.315 32.045 195.885 ;
        RECT 32.280 195.735 33.930 195.905 ;
        RECT 34.115 195.830 34.405 196.555 ;
        RECT 34.580 195.790 35.035 196.555 ;
        RECT 35.310 196.175 36.610 196.385 ;
        RECT 36.865 196.195 37.195 196.555 ;
        RECT 36.440 196.025 36.610 196.175 ;
        RECT 37.365 196.055 37.625 196.385 ;
        RECT 32.215 195.395 33.355 195.565 ;
        RECT 32.215 195.145 32.385 195.395 ;
        RECT 33.525 195.225 33.930 195.735 ;
        RECT 35.510 195.565 35.730 195.965 ;
        RECT 34.575 195.365 35.065 195.565 ;
        RECT 35.255 195.355 35.730 195.565 ;
        RECT 35.975 195.565 36.185 195.965 ;
        RECT 36.440 195.900 37.195 196.025 ;
        RECT 36.440 195.855 37.285 195.900 ;
        RECT 37.015 195.735 37.285 195.855 ;
        RECT 35.975 195.355 36.305 195.565 ;
        RECT 36.475 195.295 36.885 195.600 ;
        RECT 30.885 194.005 31.135 195.145 ;
        RECT 31.355 194.975 32.385 195.145 ;
        RECT 33.175 195.055 33.930 195.225 ;
        RECT 31.355 194.175 31.665 194.975 ;
        RECT 33.175 194.805 33.435 195.055 ;
        RECT 31.835 194.005 32.145 194.805 ;
        RECT 32.315 194.635 33.435 194.805 ;
        RECT 32.315 194.175 32.575 194.635 ;
        RECT 32.745 194.005 33.000 194.465 ;
        RECT 33.175 194.175 33.435 194.635 ;
        RECT 33.605 194.005 33.890 194.875 ;
        RECT 34.115 194.005 34.405 195.170 ;
        RECT 34.580 195.125 35.755 195.185 ;
        RECT 37.115 195.160 37.285 195.735 ;
        RECT 37.085 195.125 37.285 195.160 ;
        RECT 34.580 195.015 37.285 195.125 ;
        RECT 34.580 194.395 34.835 195.015 ;
        RECT 35.425 194.955 37.225 195.015 ;
        RECT 35.425 194.925 35.755 194.955 ;
        RECT 37.455 194.855 37.625 196.055 ;
        RECT 35.085 194.755 35.270 194.845 ;
        RECT 35.860 194.755 36.695 194.765 ;
        RECT 35.085 194.555 36.695 194.755 ;
        RECT 35.085 194.515 35.315 194.555 ;
        RECT 34.580 194.175 34.915 194.395 ;
        RECT 35.920 194.005 36.275 194.385 ;
        RECT 36.445 194.175 36.695 194.555 ;
        RECT 36.945 194.005 37.195 194.785 ;
        RECT 37.365 194.175 37.625 194.855 ;
        RECT 37.795 196.055 38.055 196.385 ;
        RECT 38.225 196.195 38.555 196.555 ;
        RECT 38.810 196.175 40.110 196.385 ;
        RECT 37.795 194.855 37.965 196.055 ;
        RECT 38.810 196.025 38.980 196.175 ;
        RECT 38.225 195.900 38.980 196.025 ;
        RECT 38.135 195.855 38.980 195.900 ;
        RECT 38.135 195.735 38.405 195.855 ;
        RECT 38.135 195.160 38.305 195.735 ;
        RECT 38.535 195.295 38.945 195.600 ;
        RECT 39.235 195.565 39.445 195.965 ;
        RECT 39.115 195.355 39.445 195.565 ;
        RECT 39.690 195.565 39.910 195.965 ;
        RECT 40.385 195.790 40.840 196.555 ;
        RECT 41.935 195.805 43.145 196.555 ;
        RECT 39.690 195.355 40.165 195.565 ;
        RECT 40.355 195.365 40.845 195.565 ;
        RECT 38.135 195.125 38.335 195.160 ;
        RECT 39.665 195.125 40.840 195.185 ;
        RECT 38.135 195.015 40.840 195.125 ;
        RECT 38.195 194.955 39.995 195.015 ;
        RECT 39.665 194.925 39.995 194.955 ;
        RECT 37.795 194.175 38.055 194.855 ;
        RECT 38.225 194.005 38.475 194.785 ;
        RECT 38.725 194.755 39.560 194.765 ;
        RECT 40.150 194.755 40.335 194.845 ;
        RECT 38.725 194.555 40.335 194.755 ;
        RECT 38.725 194.175 38.975 194.555 ;
        RECT 40.105 194.515 40.335 194.555 ;
        RECT 40.585 194.395 40.840 195.015 ;
        RECT 39.145 194.005 39.500 194.385 ;
        RECT 40.505 194.175 40.840 194.395 ;
        RECT 41.935 195.095 42.455 195.635 ;
        RECT 42.625 195.265 43.145 195.805 ;
        RECT 41.935 194.005 43.145 195.095 ;
        RECT 8.270 193.835 43.230 194.005 ;
        RECT 8.355 192.745 9.565 193.835 ;
        RECT 9.735 192.745 11.405 193.835 ;
        RECT 8.355 192.035 8.875 192.575 ;
        RECT 9.045 192.205 9.565 192.745 ;
        RECT 9.735 192.055 10.485 192.575 ;
        RECT 10.655 192.225 11.405 192.745 ;
        RECT 12.035 192.985 12.295 193.665 ;
        RECT 12.465 193.055 12.715 193.835 ;
        RECT 12.965 193.285 13.215 193.665 ;
        RECT 13.385 193.455 13.740 193.835 ;
        RECT 14.745 193.445 15.080 193.665 ;
        RECT 14.345 193.285 14.575 193.325 ;
        RECT 12.965 193.085 14.575 193.285 ;
        RECT 12.965 193.075 13.800 193.085 ;
        RECT 14.390 192.995 14.575 193.085 ;
        RECT 8.355 191.285 9.565 192.035 ;
        RECT 9.735 191.285 11.405 192.055 ;
        RECT 12.035 191.795 12.205 192.985 ;
        RECT 13.905 192.885 14.235 192.915 ;
        RECT 12.435 192.825 14.235 192.885 ;
        RECT 14.825 192.825 15.080 193.445 ;
        RECT 12.375 192.715 15.080 192.825 ;
        RECT 12.375 192.680 12.575 192.715 ;
        RECT 12.375 192.105 12.545 192.680 ;
        RECT 13.905 192.655 15.080 192.715 ;
        RECT 15.255 192.760 15.525 193.665 ;
        RECT 15.695 193.075 16.025 193.835 ;
        RECT 16.205 192.905 16.375 193.665 ;
        RECT 12.775 192.240 13.185 192.545 ;
        RECT 13.355 192.275 13.685 192.485 ;
        RECT 12.375 191.985 12.645 192.105 ;
        RECT 12.375 191.940 13.220 191.985 ;
        RECT 12.465 191.815 13.220 191.940 ;
        RECT 13.475 191.875 13.685 192.275 ;
        RECT 13.930 192.275 14.405 192.485 ;
        RECT 14.595 192.275 15.085 192.475 ;
        RECT 13.930 191.875 14.150 192.275 ;
        RECT 12.035 191.785 12.265 191.795 ;
        RECT 12.035 191.455 12.295 191.785 ;
        RECT 13.050 191.665 13.220 191.815 ;
        RECT 12.465 191.285 12.795 191.645 ;
        RECT 13.050 191.455 14.350 191.665 ;
        RECT 14.625 191.285 15.080 192.050 ;
        RECT 15.255 191.960 15.425 192.760 ;
        RECT 15.710 192.735 16.375 192.905 ;
        RECT 17.095 192.985 17.355 193.665 ;
        RECT 17.525 193.055 17.775 193.835 ;
        RECT 18.025 193.285 18.275 193.665 ;
        RECT 18.445 193.455 18.800 193.835 ;
        RECT 19.805 193.445 20.140 193.665 ;
        RECT 19.405 193.285 19.635 193.325 ;
        RECT 18.025 193.085 19.635 193.285 ;
        RECT 18.025 193.075 18.860 193.085 ;
        RECT 19.450 192.995 19.635 193.085 ;
        RECT 15.710 192.590 15.880 192.735 ;
        RECT 15.595 192.260 15.880 192.590 ;
        RECT 15.710 192.005 15.880 192.260 ;
        RECT 16.115 192.185 16.445 192.555 ;
        RECT 15.255 191.455 15.515 191.960 ;
        RECT 15.710 191.835 16.375 192.005 ;
        RECT 15.695 191.285 16.025 191.665 ;
        RECT 16.205 191.455 16.375 191.835 ;
        RECT 17.095 191.795 17.265 192.985 ;
        RECT 18.965 192.885 19.295 192.915 ;
        RECT 17.495 192.825 19.295 192.885 ;
        RECT 19.885 192.825 20.140 193.445 ;
        RECT 17.435 192.715 20.140 192.825 ;
        RECT 17.435 192.680 17.635 192.715 ;
        RECT 17.435 192.105 17.605 192.680 ;
        RECT 18.965 192.655 20.140 192.715 ;
        RECT 21.235 192.670 21.525 193.835 ;
        RECT 22.210 192.965 22.495 193.835 ;
        RECT 22.665 193.205 22.925 193.665 ;
        RECT 23.100 193.375 23.355 193.835 ;
        RECT 23.525 193.205 23.785 193.665 ;
        RECT 22.665 193.035 23.785 193.205 ;
        RECT 23.955 193.035 24.265 193.835 ;
        RECT 22.665 192.785 22.925 193.035 ;
        RECT 24.435 192.865 24.745 193.665 ;
        RECT 22.170 192.615 22.925 192.785 ;
        RECT 23.715 192.695 24.745 192.865 ;
        RECT 17.835 192.240 18.245 192.545 ;
        RECT 18.415 192.275 18.745 192.485 ;
        RECT 17.435 191.985 17.705 192.105 ;
        RECT 17.435 191.940 18.280 191.985 ;
        RECT 17.525 191.815 18.280 191.940 ;
        RECT 18.535 191.875 18.745 192.275 ;
        RECT 18.990 192.275 19.465 192.485 ;
        RECT 19.655 192.275 20.145 192.475 ;
        RECT 18.990 191.875 19.210 192.275 ;
        RECT 22.170 192.105 22.575 192.615 ;
        RECT 23.715 192.445 23.885 192.695 ;
        RECT 22.745 192.275 23.885 192.445 ;
        RECT 17.095 191.785 17.325 191.795 ;
        RECT 17.095 191.455 17.355 191.785 ;
        RECT 18.110 191.665 18.280 191.815 ;
        RECT 17.525 191.285 17.855 191.645 ;
        RECT 18.110 191.455 19.410 191.665 ;
        RECT 19.685 191.285 20.140 192.050 ;
        RECT 21.235 191.285 21.525 192.010 ;
        RECT 22.170 191.935 23.820 192.105 ;
        RECT 24.055 191.955 24.405 192.525 ;
        RECT 22.215 191.285 22.495 191.765 ;
        RECT 22.665 191.545 22.925 191.935 ;
        RECT 23.100 191.285 23.355 191.765 ;
        RECT 23.525 191.545 23.820 191.935 ;
        RECT 24.575 191.785 24.745 192.695 ;
        RECT 24.000 191.285 24.275 191.765 ;
        RECT 24.445 191.455 24.745 191.785 ;
        RECT 24.915 192.695 25.300 193.665 ;
        RECT 25.470 193.375 25.795 193.835 ;
        RECT 26.315 193.205 26.595 193.665 ;
        RECT 25.470 192.985 26.595 193.205 ;
        RECT 24.915 192.025 25.195 192.695 ;
        RECT 25.470 192.525 25.920 192.985 ;
        RECT 26.785 192.815 27.185 193.665 ;
        RECT 27.585 193.375 27.855 193.835 ;
        RECT 28.025 193.205 28.310 193.665 ;
        RECT 25.365 192.195 25.920 192.525 ;
        RECT 26.090 192.255 27.185 192.815 ;
        RECT 25.470 192.085 25.920 192.195 ;
        RECT 24.915 191.455 25.300 192.025 ;
        RECT 25.470 191.915 26.595 192.085 ;
        RECT 25.470 191.285 25.795 191.745 ;
        RECT 26.315 191.455 26.595 191.915 ;
        RECT 26.785 191.455 27.185 192.255 ;
        RECT 27.355 192.985 28.310 193.205 ;
        RECT 27.355 192.085 27.565 192.985 ;
        RECT 28.685 192.905 28.855 193.665 ;
        RECT 29.070 193.075 29.400 193.835 ;
        RECT 27.735 192.255 28.425 192.815 ;
        RECT 28.685 192.735 29.400 192.905 ;
        RECT 29.570 192.760 29.825 193.665 ;
        RECT 28.595 192.185 28.950 192.555 ;
        RECT 29.230 192.525 29.400 192.735 ;
        RECT 29.230 192.195 29.485 192.525 ;
        RECT 27.355 191.915 28.310 192.085 ;
        RECT 29.230 192.005 29.400 192.195 ;
        RECT 29.655 192.030 29.825 192.760 ;
        RECT 30.000 192.685 30.260 193.835 ;
        RECT 30.900 193.165 31.155 193.665 ;
        RECT 31.325 193.335 31.655 193.835 ;
        RECT 30.900 192.995 31.650 193.165 ;
        RECT 30.900 192.175 31.250 192.825 ;
        RECT 27.585 191.285 27.855 191.745 ;
        RECT 28.025 191.455 28.310 191.915 ;
        RECT 28.685 191.835 29.400 192.005 ;
        RECT 28.685 191.455 28.855 191.835 ;
        RECT 29.070 191.285 29.400 191.665 ;
        RECT 29.570 191.455 29.825 192.030 ;
        RECT 30.000 191.285 30.260 192.125 ;
        RECT 31.420 192.005 31.650 192.995 ;
        RECT 30.900 191.835 31.650 192.005 ;
        RECT 30.900 191.545 31.155 191.835 ;
        RECT 31.325 191.285 31.655 191.665 ;
        RECT 31.825 191.545 31.995 193.665 ;
        RECT 32.165 192.865 32.490 193.650 ;
        RECT 32.660 193.375 32.910 193.835 ;
        RECT 33.080 193.335 33.330 193.665 ;
        RECT 33.545 193.335 34.225 193.665 ;
        RECT 33.080 193.205 33.250 193.335 ;
        RECT 32.855 193.035 33.250 193.205 ;
        RECT 32.225 191.815 32.685 192.865 ;
        RECT 32.855 191.675 33.025 193.035 ;
        RECT 33.420 192.775 33.885 193.165 ;
        RECT 33.195 191.965 33.545 192.585 ;
        RECT 33.715 192.185 33.885 192.775 ;
        RECT 34.055 192.555 34.225 193.335 ;
        RECT 34.395 193.235 34.565 193.575 ;
        RECT 34.800 193.405 35.130 193.835 ;
        RECT 35.300 193.235 35.470 193.575 ;
        RECT 35.765 193.375 36.135 193.835 ;
        RECT 34.395 193.065 35.470 193.235 ;
        RECT 36.305 193.205 36.475 193.665 ;
        RECT 36.710 193.325 37.580 193.665 ;
        RECT 37.750 193.375 38.000 193.835 ;
        RECT 35.915 193.035 36.475 193.205 ;
        RECT 35.915 192.895 36.085 193.035 ;
        RECT 34.585 192.725 36.085 192.895 ;
        RECT 36.780 192.865 37.240 193.155 ;
        RECT 34.055 192.385 35.745 192.555 ;
        RECT 33.715 191.965 34.070 192.185 ;
        RECT 34.240 191.675 34.410 192.385 ;
        RECT 34.615 191.965 35.405 192.215 ;
        RECT 35.575 192.205 35.745 192.385 ;
        RECT 35.915 192.035 36.085 192.725 ;
        RECT 32.355 191.285 32.685 191.645 ;
        RECT 32.855 191.505 33.350 191.675 ;
        RECT 33.555 191.505 34.410 191.675 ;
        RECT 35.285 191.285 35.615 191.745 ;
        RECT 35.825 191.645 36.085 192.035 ;
        RECT 36.275 192.855 37.240 192.865 ;
        RECT 37.410 192.945 37.580 193.325 ;
        RECT 38.170 193.285 38.340 193.575 ;
        RECT 38.520 193.455 38.850 193.835 ;
        RECT 38.170 193.115 38.970 193.285 ;
        RECT 36.275 192.695 36.950 192.855 ;
        RECT 37.410 192.775 38.630 192.945 ;
        RECT 36.275 191.905 36.485 192.695 ;
        RECT 37.410 192.685 37.580 192.775 ;
        RECT 36.655 191.905 37.005 192.525 ;
        RECT 37.175 192.515 37.580 192.685 ;
        RECT 37.175 191.735 37.345 192.515 ;
        RECT 37.515 192.065 37.735 192.345 ;
        RECT 37.915 192.235 38.455 192.605 ;
        RECT 38.800 192.525 38.970 193.115 ;
        RECT 39.190 192.695 39.495 193.835 ;
        RECT 39.665 192.645 39.920 193.525 ;
        RECT 40.185 192.905 40.355 193.665 ;
        RECT 40.570 193.075 40.900 193.835 ;
        RECT 40.185 192.735 40.900 192.905 ;
        RECT 41.070 192.760 41.325 193.665 ;
        RECT 38.800 192.495 39.540 192.525 ;
        RECT 37.515 191.895 38.045 192.065 ;
        RECT 35.825 191.475 36.175 191.645 ;
        RECT 36.395 191.455 37.345 191.735 ;
        RECT 37.515 191.285 37.705 191.725 ;
        RECT 37.875 191.665 38.045 191.895 ;
        RECT 38.215 191.835 38.455 192.235 ;
        RECT 38.625 192.195 39.540 192.495 ;
        RECT 38.625 192.020 38.950 192.195 ;
        RECT 38.625 191.665 38.945 192.020 ;
        RECT 39.710 191.995 39.920 192.645 ;
        RECT 40.095 192.185 40.450 192.555 ;
        RECT 40.730 192.525 40.900 192.735 ;
        RECT 40.730 192.195 40.985 192.525 ;
        RECT 40.730 192.005 40.900 192.195 ;
        RECT 41.155 192.030 41.325 192.760 ;
        RECT 41.500 192.685 41.760 193.835 ;
        RECT 41.935 192.745 43.145 193.835 ;
        RECT 41.935 192.205 42.455 192.745 ;
        RECT 37.875 191.495 38.945 191.665 ;
        RECT 39.190 191.285 39.495 191.745 ;
        RECT 39.665 191.465 39.920 191.995 ;
        RECT 40.185 191.835 40.900 192.005 ;
        RECT 40.185 191.455 40.355 191.835 ;
        RECT 40.570 191.285 40.900 191.665 ;
        RECT 41.070 191.455 41.325 192.030 ;
        RECT 41.500 191.285 41.760 192.125 ;
        RECT 42.625 192.035 43.145 192.575 ;
        RECT 41.935 191.285 43.145 192.035 ;
        RECT 8.270 191.115 43.230 191.285 ;
        RECT 8.355 190.365 9.565 191.115 ;
        RECT 9.795 190.635 10.075 191.115 ;
        RECT 10.245 190.465 10.505 190.855 ;
        RECT 10.680 190.635 10.935 191.115 ;
        RECT 11.105 190.465 11.400 190.855 ;
        RECT 11.580 190.635 11.855 191.115 ;
        RECT 12.025 190.615 12.325 190.945 ;
        RECT 8.355 189.825 8.875 190.365 ;
        RECT 9.750 190.295 11.400 190.465 ;
        RECT 9.045 189.655 9.565 190.195 ;
        RECT 8.355 188.565 9.565 189.655 ;
        RECT 9.750 189.785 10.155 190.295 ;
        RECT 10.325 189.955 11.465 190.125 ;
        RECT 9.750 189.615 10.505 189.785 ;
        RECT 9.790 188.565 10.075 189.435 ;
        RECT 10.245 189.365 10.505 189.615 ;
        RECT 11.295 189.705 11.465 189.955 ;
        RECT 11.635 189.875 11.985 190.445 ;
        RECT 12.155 189.705 12.325 190.615 ;
        RECT 12.585 190.565 12.755 190.945 ;
        RECT 12.935 190.735 13.265 191.115 ;
        RECT 12.585 190.395 13.250 190.565 ;
        RECT 13.445 190.440 13.705 190.945 ;
        RECT 12.515 189.845 12.845 190.215 ;
        RECT 13.080 190.140 13.250 190.395 ;
        RECT 11.295 189.535 12.325 189.705 ;
        RECT 13.080 189.810 13.365 190.140 ;
        RECT 13.080 189.665 13.250 189.810 ;
        RECT 10.245 189.195 11.365 189.365 ;
        RECT 10.245 188.735 10.505 189.195 ;
        RECT 10.680 188.565 10.935 189.025 ;
        RECT 11.105 188.735 11.365 189.195 ;
        RECT 11.535 188.565 11.845 189.365 ;
        RECT 12.015 188.735 12.325 189.535 ;
        RECT 12.585 189.495 13.250 189.665 ;
        RECT 13.535 189.640 13.705 190.440 ;
        RECT 12.585 188.735 12.755 189.495 ;
        RECT 12.935 188.565 13.265 189.325 ;
        RECT 13.435 188.735 13.705 189.640 ;
        RECT 13.875 190.615 14.135 190.945 ;
        RECT 14.305 190.755 14.635 191.115 ;
        RECT 14.890 190.735 16.190 190.945 ;
        RECT 13.875 189.415 14.045 190.615 ;
        RECT 14.890 190.585 15.060 190.735 ;
        RECT 14.305 190.460 15.060 190.585 ;
        RECT 14.215 190.415 15.060 190.460 ;
        RECT 14.215 190.295 14.485 190.415 ;
        RECT 14.215 189.720 14.385 190.295 ;
        RECT 14.615 189.855 15.025 190.160 ;
        RECT 15.315 190.125 15.525 190.525 ;
        RECT 15.195 189.915 15.525 190.125 ;
        RECT 15.770 190.125 15.990 190.525 ;
        RECT 16.465 190.350 16.920 191.115 ;
        RECT 17.095 190.615 17.395 190.945 ;
        RECT 17.565 190.635 17.840 191.115 ;
        RECT 15.770 189.915 16.245 190.125 ;
        RECT 16.435 189.925 16.925 190.125 ;
        RECT 14.215 189.685 14.415 189.720 ;
        RECT 15.745 189.685 16.920 189.745 ;
        RECT 14.215 189.575 16.920 189.685 ;
        RECT 14.275 189.515 16.075 189.575 ;
        RECT 15.745 189.485 16.075 189.515 ;
        RECT 13.875 188.735 14.135 189.415 ;
        RECT 14.305 188.565 14.555 189.345 ;
        RECT 14.805 189.315 15.640 189.325 ;
        RECT 16.230 189.315 16.415 189.405 ;
        RECT 14.805 189.115 16.415 189.315 ;
        RECT 14.805 188.735 15.055 189.115 ;
        RECT 16.185 189.075 16.415 189.115 ;
        RECT 16.665 188.955 16.920 189.575 ;
        RECT 15.225 188.565 15.580 188.945 ;
        RECT 16.585 188.735 16.920 188.955 ;
        RECT 17.095 189.705 17.265 190.615 ;
        RECT 18.020 190.465 18.315 190.855 ;
        RECT 18.485 190.635 18.740 191.115 ;
        RECT 18.915 190.465 19.175 190.855 ;
        RECT 19.345 190.635 19.625 191.115 ;
        RECT 17.435 189.875 17.785 190.445 ;
        RECT 18.020 190.295 19.670 190.465 ;
        RECT 17.955 189.955 19.095 190.125 ;
        RECT 17.955 189.705 18.125 189.955 ;
        RECT 19.265 189.785 19.670 190.295 ;
        RECT 17.095 189.535 18.125 189.705 ;
        RECT 18.915 189.615 19.670 189.785 ;
        RECT 20.320 190.375 20.575 190.945 ;
        RECT 20.745 190.715 21.075 191.115 ;
        RECT 21.500 190.580 22.030 190.945 ;
        RECT 21.500 190.545 21.675 190.580 ;
        RECT 20.745 190.375 21.675 190.545 ;
        RECT 20.320 189.705 20.490 190.375 ;
        RECT 20.745 190.205 20.915 190.375 ;
        RECT 20.660 189.875 20.915 190.205 ;
        RECT 21.140 189.875 21.335 190.205 ;
        RECT 17.095 188.735 17.405 189.535 ;
        RECT 18.535 189.365 18.705 189.415 ;
        RECT 18.915 189.365 19.175 189.615 ;
        RECT 17.575 188.565 17.885 189.365 ;
        RECT 18.055 189.195 19.175 189.365 ;
        RECT 18.055 188.735 18.315 189.195 ;
        RECT 18.485 188.565 18.740 189.025 ;
        RECT 18.915 188.735 19.175 189.195 ;
        RECT 19.345 188.565 19.630 189.435 ;
        RECT 20.320 188.735 20.655 189.705 ;
        RECT 20.825 188.565 20.995 189.705 ;
        RECT 21.165 188.905 21.335 189.875 ;
        RECT 21.505 189.245 21.675 190.375 ;
        RECT 21.845 189.585 22.015 190.385 ;
        RECT 22.220 190.095 22.495 190.945 ;
        RECT 22.215 189.925 22.495 190.095 ;
        RECT 22.220 189.785 22.495 189.925 ;
        RECT 22.665 189.585 22.855 190.945 ;
        RECT 23.035 190.580 23.545 191.115 ;
        RECT 23.765 190.305 24.010 190.910 ;
        RECT 25.005 190.635 25.305 191.115 ;
        RECT 25.475 190.465 25.735 190.920 ;
        RECT 25.905 190.635 26.165 191.115 ;
        RECT 26.345 190.465 26.605 190.920 ;
        RECT 26.775 190.635 27.025 191.115 ;
        RECT 27.205 190.465 27.465 190.920 ;
        RECT 27.635 190.635 27.885 191.115 ;
        RECT 28.065 190.465 28.325 190.920 ;
        RECT 28.495 190.635 28.740 191.115 ;
        RECT 28.910 190.465 29.185 190.920 ;
        RECT 29.355 190.635 29.600 191.115 ;
        RECT 29.770 190.465 30.030 190.920 ;
        RECT 30.200 190.635 30.460 191.115 ;
        RECT 30.630 190.465 30.890 190.920 ;
        RECT 31.060 190.635 31.320 191.115 ;
        RECT 31.490 190.465 31.750 190.920 ;
        RECT 31.920 190.555 32.180 191.115 ;
        RECT 23.055 190.135 24.285 190.305 ;
        RECT 21.845 189.415 22.855 189.585 ;
        RECT 23.025 189.570 23.775 189.760 ;
        RECT 21.505 189.075 22.630 189.245 ;
        RECT 23.025 188.905 23.195 189.570 ;
        RECT 23.945 189.325 24.285 190.135 ;
        RECT 25.005 190.295 31.750 190.465 ;
        RECT 25.005 189.705 26.170 190.295 ;
        RECT 32.350 190.125 32.600 190.935 ;
        RECT 32.780 190.590 33.040 191.115 ;
        RECT 33.210 190.125 33.460 190.935 ;
        RECT 33.640 190.605 33.945 191.115 ;
        RECT 26.340 189.875 33.460 190.125 ;
        RECT 33.630 189.875 33.945 190.435 ;
        RECT 34.115 190.390 34.405 191.115 ;
        RECT 34.580 190.275 34.840 191.115 ;
        RECT 35.015 190.370 35.270 190.945 ;
        RECT 35.440 190.735 35.770 191.115 ;
        RECT 35.985 190.565 36.155 190.945 ;
        RECT 35.440 190.395 36.155 190.565 ;
        RECT 25.005 189.480 31.750 189.705 ;
        RECT 21.165 188.735 23.195 188.905 ;
        RECT 23.365 188.565 23.535 189.325 ;
        RECT 23.770 188.915 24.285 189.325 ;
        RECT 25.005 188.565 25.275 189.310 ;
        RECT 25.445 188.740 25.735 189.480 ;
        RECT 26.345 189.465 31.750 189.480 ;
        RECT 25.905 188.570 26.160 189.295 ;
        RECT 26.345 188.740 26.605 189.465 ;
        RECT 26.775 188.570 27.020 189.295 ;
        RECT 27.205 188.740 27.465 189.465 ;
        RECT 27.635 188.570 27.880 189.295 ;
        RECT 28.065 188.740 28.325 189.465 ;
        RECT 28.495 188.570 28.740 189.295 ;
        RECT 28.910 188.740 29.170 189.465 ;
        RECT 29.340 188.570 29.600 189.295 ;
        RECT 29.770 188.740 30.030 189.465 ;
        RECT 30.200 188.570 30.460 189.295 ;
        RECT 30.630 188.740 30.890 189.465 ;
        RECT 31.060 188.570 31.320 189.295 ;
        RECT 31.490 188.740 31.750 189.465 ;
        RECT 31.920 188.570 32.180 189.365 ;
        RECT 32.350 188.740 32.600 189.875 ;
        RECT 25.905 188.565 32.180 188.570 ;
        RECT 32.780 188.565 33.040 189.375 ;
        RECT 33.215 188.735 33.460 189.875 ;
        RECT 33.640 188.565 33.935 189.375 ;
        RECT 34.115 188.565 34.405 189.730 ;
        RECT 34.580 188.565 34.840 189.715 ;
        RECT 35.015 189.640 35.185 190.370 ;
        RECT 35.440 190.205 35.610 190.395 ;
        RECT 36.875 190.375 37.260 190.945 ;
        RECT 37.430 190.655 37.755 191.115 ;
        RECT 38.275 190.485 38.555 190.945 ;
        RECT 35.355 189.875 35.610 190.205 ;
        RECT 35.440 189.665 35.610 189.875 ;
        RECT 35.890 189.845 36.245 190.215 ;
        RECT 36.875 189.705 37.155 190.375 ;
        RECT 37.430 190.315 38.555 190.485 ;
        RECT 37.430 190.205 37.880 190.315 ;
        RECT 37.325 189.875 37.880 190.205 ;
        RECT 38.745 190.145 39.145 190.945 ;
        RECT 39.545 190.655 39.815 191.115 ;
        RECT 39.985 190.485 40.270 190.945 ;
        RECT 35.015 188.735 35.270 189.640 ;
        RECT 35.440 189.495 36.155 189.665 ;
        RECT 35.440 188.565 35.770 189.325 ;
        RECT 35.985 188.735 36.155 189.495 ;
        RECT 36.875 188.735 37.260 189.705 ;
        RECT 37.430 189.415 37.880 189.875 ;
        RECT 38.050 189.585 39.145 190.145 ;
        RECT 37.430 189.195 38.555 189.415 ;
        RECT 37.430 188.565 37.755 189.025 ;
        RECT 38.275 188.735 38.555 189.195 ;
        RECT 38.745 188.735 39.145 189.585 ;
        RECT 39.315 190.315 40.270 190.485 ;
        RECT 40.555 190.440 40.815 190.945 ;
        RECT 40.995 190.735 41.325 191.115 ;
        RECT 41.505 190.565 41.675 190.945 ;
        RECT 39.315 189.415 39.525 190.315 ;
        RECT 39.695 189.585 40.385 190.145 ;
        RECT 40.555 189.640 40.735 190.440 ;
        RECT 41.010 190.395 41.675 190.565 ;
        RECT 41.010 190.140 41.180 190.395 ;
        RECT 41.935 190.365 43.145 191.115 ;
        RECT 40.905 189.810 41.180 190.140 ;
        RECT 41.405 189.845 41.745 190.215 ;
        RECT 41.010 189.665 41.180 189.810 ;
        RECT 39.315 189.195 40.270 189.415 ;
        RECT 39.545 188.565 39.815 189.025 ;
        RECT 39.985 188.735 40.270 189.195 ;
        RECT 40.555 188.735 40.825 189.640 ;
        RECT 41.010 189.495 41.685 189.665 ;
        RECT 40.995 188.565 41.325 189.325 ;
        RECT 41.505 188.735 41.685 189.495 ;
        RECT 41.935 189.655 42.455 190.195 ;
        RECT 42.625 189.825 43.145 190.365 ;
        RECT 60.160 190.465 62.110 190.635 ;
        RECT 41.935 188.565 43.145 189.655 ;
        RECT 8.270 188.395 43.230 188.565 ;
        RECT 8.355 187.305 9.565 188.395 ;
        RECT 9.790 187.525 10.075 188.395 ;
        RECT 10.245 187.765 10.505 188.225 ;
        RECT 10.680 187.935 10.935 188.395 ;
        RECT 11.105 187.765 11.365 188.225 ;
        RECT 10.245 187.595 11.365 187.765 ;
        RECT 11.535 187.595 11.845 188.395 ;
        RECT 10.245 187.345 10.505 187.595 ;
        RECT 12.015 187.425 12.325 188.225 ;
        RECT 12.550 187.525 12.835 188.395 ;
        RECT 13.005 187.765 13.265 188.225 ;
        RECT 13.440 187.935 13.695 188.395 ;
        RECT 13.865 187.765 14.125 188.225 ;
        RECT 13.005 187.595 14.125 187.765 ;
        RECT 14.295 187.595 14.605 188.395 ;
        RECT 8.355 186.595 8.875 187.135 ;
        RECT 9.045 186.765 9.565 187.305 ;
        RECT 9.750 187.175 10.505 187.345 ;
        RECT 11.295 187.255 12.325 187.425 ;
        RECT 13.005 187.345 13.265 187.595 ;
        RECT 14.775 187.425 15.085 188.225 ;
        RECT 9.750 186.665 10.155 187.175 ;
        RECT 11.295 187.005 11.465 187.255 ;
        RECT 10.325 186.835 11.465 187.005 ;
        RECT 8.355 185.845 9.565 186.595 ;
        RECT 9.750 186.495 11.400 186.665 ;
        RECT 11.635 186.515 11.985 187.085 ;
        RECT 9.795 185.845 10.075 186.325 ;
        RECT 10.245 186.105 10.505 186.495 ;
        RECT 10.680 185.845 10.935 186.325 ;
        RECT 11.105 186.105 11.400 186.495 ;
        RECT 12.155 186.345 12.325 187.255 ;
        RECT 12.510 187.175 13.265 187.345 ;
        RECT 14.055 187.255 15.085 187.425 ;
        RECT 12.510 186.665 12.915 187.175 ;
        RECT 14.055 187.005 14.225 187.255 ;
        RECT 13.085 186.835 14.225 187.005 ;
        RECT 12.510 186.495 14.160 186.665 ;
        RECT 14.395 186.515 14.745 187.085 ;
        RECT 11.580 185.845 11.855 186.325 ;
        RECT 12.025 186.015 12.325 186.345 ;
        RECT 12.555 185.845 12.835 186.325 ;
        RECT 13.005 186.105 13.265 186.495 ;
        RECT 13.440 185.845 13.695 186.325 ;
        RECT 13.865 186.105 14.160 186.495 ;
        RECT 14.915 186.345 15.085 187.255 ;
        RECT 14.340 185.845 14.615 186.325 ;
        RECT 14.785 186.015 15.085 186.345 ;
        RECT 15.715 187.320 15.985 188.225 ;
        RECT 16.155 187.635 16.485 188.395 ;
        RECT 16.665 187.465 16.835 188.225 ;
        RECT 15.715 186.520 15.885 187.320 ;
        RECT 16.170 187.295 16.835 187.465 ;
        RECT 16.170 187.150 16.340 187.295 ;
        RECT 16.055 186.820 16.340 187.150 ;
        RECT 17.100 187.255 17.435 188.225 ;
        RECT 17.605 187.255 17.775 188.395 ;
        RECT 17.945 188.055 19.975 188.225 ;
        RECT 16.170 186.565 16.340 186.820 ;
        RECT 16.575 186.745 16.905 187.115 ;
        RECT 17.100 186.585 17.270 187.255 ;
        RECT 17.945 187.085 18.115 188.055 ;
        RECT 17.440 186.755 17.695 187.085 ;
        RECT 17.920 186.755 18.115 187.085 ;
        RECT 18.285 187.715 19.410 187.885 ;
        RECT 17.525 186.585 17.695 186.755 ;
        RECT 18.285 186.585 18.455 187.715 ;
        RECT 15.715 186.015 15.975 186.520 ;
        RECT 16.170 186.395 16.835 186.565 ;
        RECT 16.155 185.845 16.485 186.225 ;
        RECT 16.665 186.015 16.835 186.395 ;
        RECT 17.100 186.015 17.355 186.585 ;
        RECT 17.525 186.415 18.455 186.585 ;
        RECT 18.625 187.375 19.635 187.545 ;
        RECT 18.625 186.575 18.795 187.375 ;
        RECT 18.280 186.380 18.455 186.415 ;
        RECT 17.525 185.845 17.855 186.245 ;
        RECT 18.280 186.015 18.810 186.380 ;
        RECT 19.000 186.355 19.275 187.175 ;
        RECT 18.995 186.185 19.275 186.355 ;
        RECT 19.000 186.015 19.275 186.185 ;
        RECT 19.445 186.015 19.635 187.375 ;
        RECT 19.805 187.390 19.975 188.055 ;
        RECT 20.145 187.635 20.315 188.395 ;
        RECT 20.550 187.635 21.065 188.045 ;
        RECT 19.805 187.200 20.555 187.390 ;
        RECT 20.725 186.825 21.065 187.635 ;
        RECT 21.235 187.230 21.525 188.395 ;
        RECT 21.695 187.635 22.210 188.045 ;
        RECT 22.445 187.635 22.615 188.395 ;
        RECT 22.785 188.055 24.815 188.225 ;
        RECT 19.835 186.655 21.065 186.825 ;
        RECT 21.695 186.825 22.035 187.635 ;
        RECT 22.785 187.390 22.955 188.055 ;
        RECT 23.350 187.715 24.475 187.885 ;
        RECT 22.205 187.200 22.955 187.390 ;
        RECT 23.125 187.375 24.135 187.545 ;
        RECT 21.695 186.655 22.925 186.825 ;
        RECT 19.815 185.845 20.325 186.380 ;
        RECT 20.545 186.050 20.790 186.655 ;
        RECT 21.235 185.845 21.525 186.570 ;
        RECT 21.970 186.050 22.215 186.655 ;
        RECT 22.435 185.845 22.945 186.380 ;
        RECT 23.125 186.015 23.315 187.375 ;
        RECT 23.485 187.035 23.760 187.175 ;
        RECT 23.485 186.865 23.765 187.035 ;
        RECT 23.485 186.015 23.760 186.865 ;
        RECT 23.965 186.575 24.135 187.375 ;
        RECT 24.305 186.585 24.475 187.715 ;
        RECT 24.645 187.085 24.815 188.055 ;
        RECT 24.985 187.255 25.155 188.395 ;
        RECT 25.325 187.255 25.660 188.225 ;
        RECT 24.645 186.755 24.840 187.085 ;
        RECT 25.065 186.755 25.320 187.085 ;
        RECT 25.065 186.585 25.235 186.755 ;
        RECT 25.490 186.585 25.660 187.255 ;
        RECT 24.305 186.415 25.235 186.585 ;
        RECT 24.305 186.380 24.480 186.415 ;
        RECT 23.950 186.015 24.480 186.380 ;
        RECT 24.905 185.845 25.235 186.245 ;
        RECT 25.405 186.015 25.660 186.585 ;
        RECT 26.295 187.425 26.605 188.225 ;
        RECT 26.775 187.595 27.085 188.395 ;
        RECT 27.255 187.765 27.515 188.225 ;
        RECT 27.685 187.935 27.940 188.395 ;
        RECT 28.115 187.765 28.375 188.225 ;
        RECT 27.255 187.595 28.375 187.765 ;
        RECT 26.295 187.255 27.325 187.425 ;
        RECT 26.295 186.345 26.465 187.255 ;
        RECT 26.635 186.515 26.985 187.085 ;
        RECT 27.155 187.005 27.325 187.255 ;
        RECT 28.115 187.345 28.375 187.595 ;
        RECT 28.545 187.525 28.830 188.395 ;
        RECT 29.065 187.585 29.360 188.395 ;
        RECT 28.115 187.175 28.870 187.345 ;
        RECT 27.155 186.835 28.295 187.005 ;
        RECT 28.465 186.665 28.870 187.175 ;
        RECT 29.540 187.085 29.785 188.225 ;
        RECT 29.960 187.585 30.220 188.395 ;
        RECT 30.820 188.390 37.095 188.395 ;
        RECT 30.400 187.085 30.650 188.220 ;
        RECT 30.820 187.595 31.080 188.390 ;
        RECT 31.250 187.495 31.510 188.220 ;
        RECT 31.680 187.665 31.940 188.390 ;
        RECT 32.110 187.495 32.370 188.220 ;
        RECT 32.540 187.665 32.800 188.390 ;
        RECT 32.970 187.495 33.230 188.220 ;
        RECT 33.400 187.665 33.660 188.390 ;
        RECT 33.830 187.495 34.090 188.220 ;
        RECT 34.260 187.665 34.505 188.390 ;
        RECT 34.675 187.495 34.935 188.220 ;
        RECT 35.120 187.665 35.365 188.390 ;
        RECT 35.535 187.495 35.795 188.220 ;
        RECT 35.980 187.665 36.225 188.390 ;
        RECT 36.395 187.495 36.655 188.220 ;
        RECT 36.840 187.665 37.095 188.390 ;
        RECT 31.250 187.480 36.655 187.495 ;
        RECT 37.265 187.480 37.555 188.220 ;
        RECT 37.725 187.650 37.995 188.395 ;
        RECT 31.250 187.255 37.995 187.480 ;
        RECT 27.220 186.495 28.870 186.665 ;
        RECT 29.055 186.525 29.370 187.085 ;
        RECT 29.540 186.835 36.660 187.085 ;
        RECT 26.295 186.015 26.595 186.345 ;
        RECT 26.765 185.845 27.040 186.325 ;
        RECT 27.220 186.105 27.515 186.495 ;
        RECT 27.685 185.845 27.940 186.325 ;
        RECT 28.115 186.105 28.375 186.495 ;
        RECT 28.545 185.845 28.825 186.325 ;
        RECT 29.055 185.845 29.360 186.355 ;
        RECT 29.540 186.025 29.790 186.835 ;
        RECT 29.960 185.845 30.220 186.370 ;
        RECT 30.400 186.025 30.650 186.835 ;
        RECT 36.830 186.665 37.995 187.255 ;
        RECT 31.250 186.495 37.995 186.665 ;
        RECT 38.255 187.255 38.640 188.225 ;
        RECT 38.810 187.935 39.135 188.395 ;
        RECT 39.655 187.765 39.935 188.225 ;
        RECT 38.810 187.545 39.935 187.765 ;
        RECT 38.255 186.585 38.535 187.255 ;
        RECT 38.810 187.085 39.260 187.545 ;
        RECT 40.125 187.375 40.525 188.225 ;
        RECT 40.925 187.935 41.195 188.395 ;
        RECT 41.365 187.765 41.650 188.225 ;
        RECT 38.705 186.755 39.260 187.085 ;
        RECT 39.430 186.815 40.525 187.375 ;
        RECT 38.810 186.645 39.260 186.755 ;
        RECT 30.820 185.845 31.080 186.405 ;
        RECT 31.250 186.040 31.510 186.495 ;
        RECT 31.680 185.845 31.940 186.325 ;
        RECT 32.110 186.040 32.370 186.495 ;
        RECT 32.540 185.845 32.800 186.325 ;
        RECT 32.970 186.040 33.230 186.495 ;
        RECT 33.400 185.845 33.645 186.325 ;
        RECT 33.815 186.040 34.090 186.495 ;
        RECT 34.260 185.845 34.505 186.325 ;
        RECT 34.675 186.040 34.935 186.495 ;
        RECT 35.115 185.845 35.365 186.325 ;
        RECT 35.535 186.040 35.795 186.495 ;
        RECT 35.975 185.845 36.225 186.325 ;
        RECT 36.395 186.040 36.655 186.495 ;
        RECT 36.835 185.845 37.095 186.325 ;
        RECT 37.265 186.040 37.525 186.495 ;
        RECT 37.695 185.845 37.995 186.325 ;
        RECT 38.255 186.015 38.640 186.585 ;
        RECT 38.810 186.475 39.935 186.645 ;
        RECT 38.810 185.845 39.135 186.305 ;
        RECT 39.655 186.015 39.935 186.475 ;
        RECT 40.125 186.015 40.525 186.815 ;
        RECT 40.695 187.545 41.650 187.765 ;
        RECT 40.695 186.645 40.905 187.545 ;
        RECT 41.075 186.815 41.765 187.375 ;
        RECT 41.935 187.305 43.145 188.395 ;
        RECT 60.160 188.130 60.330 190.465 ;
        RECT 60.960 189.955 61.310 190.125 ;
        RECT 58.510 187.960 60.335 188.130 ;
        RECT 41.935 186.765 42.455 187.305 ;
        RECT 40.695 186.475 41.650 186.645 ;
        RECT 42.625 186.595 43.145 187.135 ;
        RECT 58.850 186.820 59.060 187.960 ;
        RECT 59.730 187.955 60.335 187.960 ;
        RECT 59.230 186.870 59.560 187.790 ;
        RECT 60.160 186.975 60.330 187.955 ;
        RECT 60.730 187.700 60.900 189.740 ;
        RECT 61.370 187.700 61.540 189.740 ;
        RECT 60.960 187.315 61.310 187.485 ;
        RECT 61.940 186.975 62.110 190.465 ;
        RECT 59.230 186.810 59.975 186.870 ;
        RECT 59.330 186.700 59.975 186.810 ;
        RECT 60.160 186.805 62.110 186.975 ;
        RECT 40.925 185.845 41.195 186.305 ;
        RECT 41.365 186.015 41.650 186.475 ;
        RECT 41.935 185.845 43.145 186.595 ;
        RECT 58.830 186.585 59.160 186.640 ;
        RECT 58.370 186.405 59.160 186.585 ;
        RECT 58.830 186.400 59.160 186.405 ;
        RECT 8.270 185.675 43.230 185.845 ;
        RECT 8.355 184.925 9.565 185.675 ;
        RECT 8.355 184.385 8.875 184.925 ;
        RECT 9.735 184.905 11.405 185.675 ;
        RECT 12.055 184.945 12.345 185.675 ;
        RECT 9.045 184.215 9.565 184.755 ;
        RECT 9.735 184.385 10.485 184.905 ;
        RECT 10.655 184.215 11.405 184.735 ;
        RECT 12.045 184.435 12.345 184.765 ;
        RECT 12.525 184.745 12.755 185.385 ;
        RECT 12.935 185.125 13.245 185.495 ;
        RECT 13.425 185.305 14.095 185.675 ;
        RECT 12.935 184.925 14.165 185.125 ;
        RECT 12.525 184.435 13.050 184.745 ;
        RECT 13.230 184.435 13.695 184.745 ;
        RECT 13.875 184.255 14.165 184.925 ;
        RECT 8.355 183.125 9.565 184.215 ;
        RECT 9.735 183.125 11.405 184.215 ;
        RECT 12.055 184.015 13.215 184.255 ;
        RECT 12.055 183.305 12.315 184.015 ;
        RECT 12.485 183.125 12.815 183.835 ;
        RECT 12.985 183.305 13.215 184.015 ;
        RECT 13.395 184.035 14.165 184.255 ;
        RECT 13.395 183.305 13.665 184.035 ;
        RECT 13.845 183.125 14.185 183.855 ;
        RECT 14.355 183.305 14.615 185.495 ;
        RECT 14.885 185.125 15.055 185.415 ;
        RECT 15.225 185.295 15.555 185.675 ;
        RECT 14.885 184.955 15.550 185.125 ;
        RECT 14.800 184.135 15.150 184.785 ;
        RECT 15.320 183.965 15.550 184.955 ;
        RECT 14.885 183.795 15.550 183.965 ;
        RECT 14.885 183.295 15.055 183.795 ;
        RECT 15.225 183.125 15.555 183.625 ;
        RECT 15.725 183.295 15.950 185.415 ;
        RECT 16.165 185.295 16.495 185.675 ;
        RECT 16.665 185.125 16.835 185.455 ;
        RECT 17.135 185.295 18.150 185.495 ;
        RECT 16.140 184.935 16.835 185.125 ;
        RECT 16.140 183.965 16.310 184.935 ;
        RECT 16.480 184.135 16.890 184.755 ;
        RECT 17.060 184.185 17.280 185.055 ;
        RECT 17.460 184.745 17.810 185.115 ;
        RECT 17.980 184.565 18.150 185.295 ;
        RECT 18.320 185.235 18.730 185.675 ;
        RECT 19.020 185.035 19.270 185.465 ;
        RECT 19.470 185.215 19.790 185.675 ;
        RECT 20.350 185.285 21.200 185.455 ;
        RECT 18.320 184.695 18.730 185.025 ;
        RECT 19.020 184.695 19.440 185.035 ;
        RECT 17.730 184.525 18.150 184.565 ;
        RECT 17.730 184.355 19.080 184.525 ;
        RECT 16.140 183.795 16.835 183.965 ;
        RECT 17.060 183.805 17.560 184.185 ;
        RECT 16.165 183.125 16.495 183.625 ;
        RECT 16.665 183.295 16.835 183.795 ;
        RECT 17.730 183.510 17.900 184.355 ;
        RECT 18.830 184.195 19.080 184.355 ;
        RECT 18.070 183.925 18.320 184.185 ;
        RECT 19.250 183.925 19.440 184.695 ;
        RECT 18.070 183.675 19.440 183.925 ;
        RECT 19.610 184.865 20.860 185.035 ;
        RECT 19.610 184.105 19.780 184.865 ;
        RECT 20.530 184.745 20.860 184.865 ;
        RECT 19.950 184.285 20.130 184.695 ;
        RECT 21.030 184.525 21.200 185.285 ;
        RECT 21.400 185.195 22.060 185.675 ;
        RECT 22.240 185.080 22.560 185.410 ;
        RECT 21.390 184.755 22.050 185.025 ;
        RECT 21.390 184.695 21.720 184.755 ;
        RECT 21.870 184.525 22.200 184.585 ;
        RECT 20.300 184.355 22.200 184.525 ;
        RECT 19.610 183.795 20.130 184.105 ;
        RECT 20.300 183.845 20.470 184.355 ;
        RECT 22.370 184.185 22.560 185.080 ;
        RECT 20.640 184.015 22.560 184.185 ;
        RECT 22.240 183.995 22.560 184.015 ;
        RECT 22.760 184.765 23.010 185.415 ;
        RECT 23.190 185.215 23.475 185.675 ;
        RECT 23.655 184.965 23.910 185.495 ;
        RECT 22.760 184.435 23.560 184.765 ;
        RECT 20.300 183.675 21.510 183.845 ;
        RECT 17.070 183.340 17.900 183.510 ;
        RECT 18.140 183.125 18.520 183.505 ;
        RECT 18.700 183.385 18.870 183.675 ;
        RECT 20.300 183.595 20.470 183.675 ;
        RECT 19.040 183.125 19.370 183.505 ;
        RECT 19.840 183.345 20.470 183.595 ;
        RECT 20.650 183.125 21.070 183.505 ;
        RECT 21.270 183.385 21.510 183.675 ;
        RECT 21.740 183.125 22.070 183.815 ;
        RECT 22.240 183.385 22.410 183.995 ;
        RECT 22.760 183.845 23.010 184.435 ;
        RECT 23.730 184.105 23.910 184.965 ;
        RECT 24.460 185.125 24.715 185.415 ;
        RECT 24.885 185.295 25.215 185.675 ;
        RECT 24.460 184.955 25.210 185.125 ;
        RECT 24.460 184.135 24.810 184.785 ;
        RECT 22.680 183.335 23.010 183.845 ;
        RECT 23.190 183.125 23.475 183.925 ;
        RECT 23.655 183.635 23.910 184.105 ;
        RECT 24.980 183.965 25.210 184.955 ;
        RECT 24.460 183.795 25.210 183.965 ;
        RECT 23.655 183.465 23.995 183.635 ;
        RECT 23.655 183.435 23.910 183.465 ;
        RECT 24.460 183.295 24.715 183.795 ;
        RECT 24.885 183.125 25.215 183.625 ;
        RECT 25.385 183.295 25.555 185.415 ;
        RECT 25.915 185.315 26.245 185.675 ;
        RECT 26.415 185.285 26.910 185.455 ;
        RECT 27.115 185.285 27.970 185.455 ;
        RECT 25.785 184.095 26.245 185.145 ;
        RECT 25.725 183.310 26.050 184.095 ;
        RECT 26.415 183.925 26.585 185.285 ;
        RECT 26.755 184.375 27.105 184.995 ;
        RECT 27.275 184.775 27.630 184.995 ;
        RECT 27.275 184.185 27.445 184.775 ;
        RECT 27.800 184.575 27.970 185.285 ;
        RECT 28.845 185.215 29.175 185.675 ;
        RECT 29.385 185.315 29.735 185.485 ;
        RECT 28.175 184.745 28.965 184.995 ;
        RECT 29.385 184.925 29.645 185.315 ;
        RECT 29.955 185.225 30.905 185.505 ;
        RECT 31.075 185.235 31.265 185.675 ;
        RECT 31.435 185.295 32.505 185.465 ;
        RECT 29.135 184.575 29.305 184.755 ;
        RECT 26.415 183.755 26.810 183.925 ;
        RECT 26.980 183.795 27.445 184.185 ;
        RECT 27.615 184.405 29.305 184.575 ;
        RECT 26.640 183.625 26.810 183.755 ;
        RECT 27.615 183.625 27.785 184.405 ;
        RECT 29.475 184.235 29.645 184.925 ;
        RECT 28.145 184.065 29.645 184.235 ;
        RECT 29.835 184.265 30.045 185.055 ;
        RECT 30.215 184.435 30.565 185.055 ;
        RECT 30.735 184.445 30.905 185.225 ;
        RECT 31.435 185.065 31.605 185.295 ;
        RECT 31.075 184.895 31.605 185.065 ;
        RECT 31.075 184.615 31.295 184.895 ;
        RECT 31.775 184.725 32.015 185.125 ;
        RECT 30.735 184.275 31.140 184.445 ;
        RECT 31.475 184.355 32.015 184.725 ;
        RECT 32.185 184.940 32.505 185.295 ;
        RECT 32.750 185.215 33.055 185.675 ;
        RECT 33.225 184.965 33.480 185.495 ;
        RECT 32.185 184.765 32.510 184.940 ;
        RECT 32.185 184.465 33.100 184.765 ;
        RECT 32.360 184.435 33.100 184.465 ;
        RECT 29.835 184.105 30.510 184.265 ;
        RECT 30.970 184.185 31.140 184.275 ;
        RECT 29.835 184.095 30.800 184.105 ;
        RECT 29.475 183.925 29.645 184.065 ;
        RECT 26.220 183.125 26.470 183.585 ;
        RECT 26.640 183.295 26.890 183.625 ;
        RECT 27.105 183.295 27.785 183.625 ;
        RECT 27.955 183.725 29.030 183.895 ;
        RECT 29.475 183.755 30.035 183.925 ;
        RECT 30.340 183.805 30.800 184.095 ;
        RECT 30.970 184.015 32.190 184.185 ;
        RECT 27.955 183.385 28.125 183.725 ;
        RECT 28.360 183.125 28.690 183.555 ;
        RECT 28.860 183.385 29.030 183.725 ;
        RECT 29.325 183.125 29.695 183.585 ;
        RECT 29.865 183.295 30.035 183.755 ;
        RECT 30.970 183.635 31.140 184.015 ;
        RECT 32.360 183.845 32.530 184.435 ;
        RECT 33.270 184.315 33.480 184.965 ;
        RECT 34.115 184.950 34.405 185.675 ;
        RECT 30.270 183.295 31.140 183.635 ;
        RECT 31.730 183.675 32.530 183.845 ;
        RECT 31.310 183.125 31.560 183.585 ;
        RECT 31.730 183.385 31.900 183.675 ;
        RECT 32.080 183.125 32.410 183.505 ;
        RECT 32.750 183.125 33.055 184.265 ;
        RECT 33.225 183.435 33.480 184.315 ;
        RECT 34.575 184.935 34.960 185.505 ;
        RECT 35.130 185.215 35.455 185.675 ;
        RECT 35.975 185.045 36.255 185.505 ;
        RECT 34.115 183.125 34.405 184.290 ;
        RECT 34.575 184.265 34.855 184.935 ;
        RECT 35.130 184.875 36.255 185.045 ;
        RECT 35.130 184.765 35.580 184.875 ;
        RECT 35.025 184.435 35.580 184.765 ;
        RECT 36.445 184.705 36.845 185.505 ;
        RECT 37.245 185.215 37.515 185.675 ;
        RECT 37.685 185.045 37.970 185.505 ;
        RECT 34.575 183.295 34.960 184.265 ;
        RECT 35.130 183.975 35.580 184.435 ;
        RECT 35.750 184.145 36.845 184.705 ;
        RECT 35.130 183.755 36.255 183.975 ;
        RECT 35.130 183.125 35.455 183.585 ;
        RECT 35.975 183.295 36.255 183.755 ;
        RECT 36.445 183.295 36.845 184.145 ;
        RECT 37.015 184.875 37.970 185.045 ;
        RECT 38.720 184.910 39.175 185.675 ;
        RECT 39.450 185.295 40.750 185.505 ;
        RECT 41.005 185.315 41.335 185.675 ;
        RECT 40.580 185.145 40.750 185.295 ;
        RECT 41.505 185.175 41.765 185.505 ;
        RECT 41.535 185.165 41.765 185.175 ;
        RECT 37.015 183.975 37.225 184.875 ;
        RECT 37.395 184.145 38.085 184.705 ;
        RECT 39.650 184.685 39.870 185.085 ;
        RECT 38.715 184.485 39.205 184.685 ;
        RECT 39.395 184.475 39.870 184.685 ;
        RECT 40.115 184.685 40.325 185.085 ;
        RECT 40.580 185.020 41.335 185.145 ;
        RECT 40.580 184.975 41.425 185.020 ;
        RECT 41.155 184.855 41.425 184.975 ;
        RECT 40.115 184.475 40.445 184.685 ;
        RECT 40.615 184.415 41.025 184.720 ;
        RECT 38.720 184.245 39.895 184.305 ;
        RECT 41.255 184.280 41.425 184.855 ;
        RECT 41.225 184.245 41.425 184.280 ;
        RECT 38.720 184.135 41.425 184.245 ;
        RECT 37.015 183.755 37.970 183.975 ;
        RECT 37.245 183.125 37.515 183.585 ;
        RECT 37.685 183.295 37.970 183.755 ;
        RECT 38.720 183.515 38.975 184.135 ;
        RECT 39.565 184.075 41.365 184.135 ;
        RECT 39.565 184.045 39.895 184.075 ;
        RECT 41.595 183.975 41.765 185.165 ;
        RECT 41.935 184.925 43.145 185.675 ;
        RECT 58.830 185.410 59.060 186.230 ;
        RECT 59.330 186.210 59.560 186.700 ;
        RECT 59.230 185.580 59.560 186.210 ;
        RECT 60.270 186.205 62.020 186.375 ;
        RECT 60.270 185.425 60.440 186.205 ;
        RECT 60.980 185.695 61.310 185.865 ;
        RECT 59.730 185.410 60.445 185.425 ;
        RECT 58.510 185.250 60.445 185.410 ;
        RECT 58.510 185.240 59.890 185.250 ;
        RECT 39.225 183.875 39.410 183.965 ;
        RECT 40.000 183.875 40.835 183.885 ;
        RECT 39.225 183.675 40.835 183.875 ;
        RECT 39.225 183.635 39.455 183.675 ;
        RECT 38.720 183.295 39.055 183.515 ;
        RECT 40.060 183.125 40.415 183.505 ;
        RECT 40.585 183.295 40.835 183.675 ;
        RECT 41.085 183.125 41.335 183.905 ;
        RECT 41.505 183.295 41.765 183.975 ;
        RECT 41.935 184.215 42.455 184.755 ;
        RECT 42.625 184.385 43.145 184.925 ;
        RECT 60.270 184.385 60.440 185.250 ;
        RECT 60.840 185.065 61.010 185.525 ;
        RECT 61.280 185.065 61.450 185.525 ;
        RECT 60.980 184.725 61.310 184.895 ;
        RECT 61.850 184.385 62.020 186.205 ;
        RECT 60.270 184.215 62.020 184.385 ;
        RECT 41.935 183.125 43.145 184.215 ;
        RECT 8.270 182.955 43.230 183.125 ;
        RECT 8.355 181.865 9.565 182.955 ;
        RECT 9.735 181.865 11.405 182.955 ;
        RECT 12.040 182.285 12.295 182.785 ;
        RECT 12.465 182.455 12.795 182.955 ;
        RECT 12.040 182.115 12.790 182.285 ;
        RECT 8.355 181.155 8.875 181.695 ;
        RECT 9.045 181.325 9.565 181.865 ;
        RECT 9.735 181.175 10.485 181.695 ;
        RECT 10.655 181.345 11.405 181.865 ;
        RECT 12.040 181.295 12.390 181.945 ;
        RECT 8.355 180.405 9.565 181.155 ;
        RECT 9.735 180.405 11.405 181.175 ;
        RECT 12.560 181.125 12.790 182.115 ;
        RECT 12.040 180.955 12.790 181.125 ;
        RECT 12.040 180.665 12.295 180.955 ;
        RECT 12.465 180.405 12.795 180.785 ;
        RECT 12.965 180.665 13.135 182.785 ;
        RECT 13.305 181.985 13.630 182.770 ;
        RECT 13.800 182.495 14.050 182.955 ;
        RECT 14.220 182.455 14.470 182.785 ;
        RECT 14.685 182.455 15.365 182.785 ;
        RECT 14.220 182.325 14.390 182.455 ;
        RECT 13.995 182.155 14.390 182.325 ;
        RECT 13.365 180.935 13.825 181.985 ;
        RECT 13.995 180.795 14.165 182.155 ;
        RECT 14.560 181.895 15.025 182.285 ;
        RECT 14.335 181.085 14.685 181.705 ;
        RECT 14.855 181.305 15.025 181.895 ;
        RECT 15.195 181.675 15.365 182.455 ;
        RECT 15.535 182.355 15.705 182.695 ;
        RECT 15.940 182.525 16.270 182.955 ;
        RECT 16.440 182.355 16.610 182.695 ;
        RECT 16.905 182.495 17.275 182.955 ;
        RECT 15.535 182.185 16.610 182.355 ;
        RECT 17.445 182.325 17.615 182.785 ;
        RECT 17.850 182.445 18.720 182.785 ;
        RECT 18.890 182.495 19.140 182.955 ;
        RECT 17.055 182.155 17.615 182.325 ;
        RECT 17.055 182.015 17.225 182.155 ;
        RECT 15.725 181.845 17.225 182.015 ;
        RECT 17.920 181.985 18.380 182.275 ;
        RECT 15.195 181.505 16.885 181.675 ;
        RECT 14.855 181.085 15.210 181.305 ;
        RECT 15.380 180.795 15.550 181.505 ;
        RECT 15.755 181.085 16.545 181.335 ;
        RECT 16.715 181.325 16.885 181.505 ;
        RECT 17.055 181.155 17.225 181.845 ;
        RECT 13.495 180.405 13.825 180.765 ;
        RECT 13.995 180.625 14.490 180.795 ;
        RECT 14.695 180.625 15.550 180.795 ;
        RECT 16.425 180.405 16.755 180.865 ;
        RECT 16.965 180.765 17.225 181.155 ;
        RECT 17.415 181.975 18.380 181.985 ;
        RECT 18.550 182.065 18.720 182.445 ;
        RECT 19.310 182.405 19.480 182.695 ;
        RECT 19.660 182.575 19.990 182.955 ;
        RECT 19.310 182.235 20.110 182.405 ;
        RECT 17.415 181.815 18.090 181.975 ;
        RECT 18.550 181.895 19.770 182.065 ;
        RECT 17.415 181.025 17.625 181.815 ;
        RECT 18.550 181.805 18.720 181.895 ;
        RECT 17.795 181.025 18.145 181.645 ;
        RECT 18.315 181.635 18.720 181.805 ;
        RECT 18.315 180.855 18.485 181.635 ;
        RECT 18.655 181.185 18.875 181.465 ;
        RECT 19.055 181.355 19.595 181.725 ;
        RECT 19.940 181.645 20.110 182.235 ;
        RECT 20.330 181.815 20.635 182.955 ;
        RECT 20.805 181.765 21.060 182.645 ;
        RECT 21.235 181.790 21.525 182.955 ;
        RECT 21.785 182.025 21.955 182.785 ;
        RECT 22.135 182.195 22.465 182.955 ;
        RECT 21.785 181.855 22.450 182.025 ;
        RECT 22.635 181.880 22.905 182.785 ;
        RECT 19.940 181.615 20.680 181.645 ;
        RECT 18.655 181.015 19.185 181.185 ;
        RECT 16.965 180.595 17.315 180.765 ;
        RECT 17.535 180.575 18.485 180.855 ;
        RECT 18.655 180.405 18.845 180.845 ;
        RECT 19.015 180.785 19.185 181.015 ;
        RECT 19.355 180.955 19.595 181.355 ;
        RECT 19.765 181.315 20.680 181.615 ;
        RECT 19.765 181.140 20.090 181.315 ;
        RECT 19.765 180.785 20.085 181.140 ;
        RECT 20.850 181.115 21.060 181.765 ;
        RECT 22.280 181.710 22.450 181.855 ;
        RECT 21.715 181.305 22.045 181.675 ;
        RECT 22.280 181.380 22.565 181.710 ;
        RECT 19.015 180.615 20.085 180.785 ;
        RECT 20.330 180.405 20.635 180.865 ;
        RECT 20.805 180.585 21.060 181.115 ;
        RECT 21.235 180.405 21.525 181.130 ;
        RECT 22.280 181.125 22.450 181.380 ;
        RECT 21.785 180.955 22.450 181.125 ;
        RECT 22.735 181.080 22.905 181.880 ;
        RECT 21.785 180.575 21.955 180.955 ;
        RECT 22.135 180.405 22.465 180.785 ;
        RECT 22.645 180.575 22.905 181.080 ;
        RECT 23.080 181.765 23.335 182.645 ;
        RECT 23.505 181.815 23.810 182.955 ;
        RECT 24.150 182.575 24.480 182.955 ;
        RECT 24.660 182.405 24.830 182.695 ;
        RECT 25.000 182.495 25.250 182.955 ;
        RECT 24.030 182.235 24.830 182.405 ;
        RECT 25.420 182.445 26.290 182.785 ;
        RECT 23.080 181.115 23.290 181.765 ;
        RECT 24.030 181.645 24.200 182.235 ;
        RECT 25.420 182.065 25.590 182.445 ;
        RECT 26.525 182.325 26.695 182.785 ;
        RECT 26.865 182.495 27.235 182.955 ;
        RECT 27.530 182.355 27.700 182.695 ;
        RECT 27.870 182.525 28.200 182.955 ;
        RECT 28.435 182.355 28.605 182.695 ;
        RECT 24.370 181.895 25.590 182.065 ;
        RECT 25.760 181.985 26.220 182.275 ;
        RECT 26.525 182.155 27.085 182.325 ;
        RECT 27.530 182.185 28.605 182.355 ;
        RECT 28.775 182.455 29.455 182.785 ;
        RECT 29.670 182.455 29.920 182.785 ;
        RECT 30.090 182.495 30.340 182.955 ;
        RECT 26.915 182.015 27.085 182.155 ;
        RECT 25.760 181.975 26.725 181.985 ;
        RECT 25.420 181.805 25.590 181.895 ;
        RECT 26.050 181.815 26.725 181.975 ;
        RECT 23.460 181.615 24.200 181.645 ;
        RECT 23.460 181.315 24.375 181.615 ;
        RECT 24.050 181.140 24.375 181.315 ;
        RECT 23.080 180.585 23.335 181.115 ;
        RECT 23.505 180.405 23.810 180.865 ;
        RECT 24.055 180.785 24.375 181.140 ;
        RECT 24.545 181.355 25.085 181.725 ;
        RECT 25.420 181.635 25.825 181.805 ;
        RECT 24.545 180.955 24.785 181.355 ;
        RECT 25.265 181.185 25.485 181.465 ;
        RECT 24.955 181.015 25.485 181.185 ;
        RECT 24.955 180.785 25.125 181.015 ;
        RECT 25.655 180.855 25.825 181.635 ;
        RECT 25.995 181.025 26.345 181.645 ;
        RECT 26.515 181.025 26.725 181.815 ;
        RECT 26.915 181.845 28.415 182.015 ;
        RECT 26.915 181.155 27.085 181.845 ;
        RECT 28.775 181.675 28.945 182.455 ;
        RECT 29.750 182.325 29.920 182.455 ;
        RECT 27.255 181.505 28.945 181.675 ;
        RECT 29.115 181.895 29.580 182.285 ;
        RECT 29.750 182.155 30.145 182.325 ;
        RECT 27.255 181.325 27.425 181.505 ;
        RECT 24.055 180.615 25.125 180.785 ;
        RECT 25.295 180.405 25.485 180.845 ;
        RECT 25.655 180.575 26.605 180.855 ;
        RECT 26.915 180.765 27.175 181.155 ;
        RECT 27.595 181.085 28.385 181.335 ;
        RECT 26.825 180.595 27.175 180.765 ;
        RECT 27.385 180.405 27.715 180.865 ;
        RECT 28.590 180.795 28.760 181.505 ;
        RECT 29.115 181.305 29.285 181.895 ;
        RECT 28.930 181.085 29.285 181.305 ;
        RECT 29.455 181.085 29.805 181.705 ;
        RECT 29.975 180.795 30.145 182.155 ;
        RECT 30.510 181.985 30.835 182.770 ;
        RECT 30.315 180.935 30.775 181.985 ;
        RECT 28.590 180.625 29.445 180.795 ;
        RECT 29.650 180.625 30.145 180.795 ;
        RECT 30.315 180.405 30.645 180.765 ;
        RECT 31.005 180.665 31.175 182.785 ;
        RECT 31.345 182.455 31.675 182.955 ;
        RECT 31.845 182.285 32.100 182.785 ;
        RECT 31.350 182.115 32.100 182.285 ;
        RECT 32.280 182.285 32.535 182.785 ;
        RECT 32.705 182.455 33.035 182.955 ;
        RECT 32.280 182.115 33.030 182.285 ;
        RECT 31.350 181.125 31.580 182.115 ;
        RECT 31.750 181.295 32.100 181.945 ;
        RECT 32.280 181.295 32.630 181.945 ;
        RECT 32.800 181.125 33.030 182.115 ;
        RECT 31.350 180.955 32.100 181.125 ;
        RECT 31.345 180.405 31.675 180.785 ;
        RECT 31.845 180.665 32.100 180.955 ;
        RECT 32.280 180.955 33.030 181.125 ;
        RECT 32.280 180.665 32.535 180.955 ;
        RECT 32.705 180.405 33.035 180.785 ;
        RECT 33.205 180.665 33.375 182.785 ;
        RECT 33.545 181.985 33.870 182.770 ;
        RECT 34.040 182.495 34.290 182.955 ;
        RECT 34.460 182.455 34.710 182.785 ;
        RECT 34.925 182.455 35.605 182.785 ;
        RECT 34.460 182.325 34.630 182.455 ;
        RECT 34.235 182.155 34.630 182.325 ;
        RECT 33.605 180.935 34.065 181.985 ;
        RECT 34.235 180.795 34.405 182.155 ;
        RECT 34.800 181.895 35.265 182.285 ;
        RECT 34.575 181.085 34.925 181.705 ;
        RECT 35.095 181.305 35.265 181.895 ;
        RECT 35.435 181.675 35.605 182.455 ;
        RECT 35.775 182.355 35.945 182.695 ;
        RECT 36.180 182.525 36.510 182.955 ;
        RECT 36.680 182.355 36.850 182.695 ;
        RECT 37.145 182.495 37.515 182.955 ;
        RECT 35.775 182.185 36.850 182.355 ;
        RECT 37.685 182.325 37.855 182.785 ;
        RECT 38.090 182.445 38.960 182.785 ;
        RECT 39.130 182.495 39.380 182.955 ;
        RECT 37.295 182.155 37.855 182.325 ;
        RECT 37.295 182.015 37.465 182.155 ;
        RECT 35.965 181.845 37.465 182.015 ;
        RECT 38.160 181.985 38.620 182.275 ;
        RECT 35.435 181.505 37.125 181.675 ;
        RECT 35.095 181.085 35.450 181.305 ;
        RECT 35.620 180.795 35.790 181.505 ;
        RECT 35.995 181.085 36.785 181.335 ;
        RECT 36.955 181.325 37.125 181.505 ;
        RECT 37.295 181.155 37.465 181.845 ;
        RECT 33.735 180.405 34.065 180.765 ;
        RECT 34.235 180.625 34.730 180.795 ;
        RECT 34.935 180.625 35.790 180.795 ;
        RECT 36.665 180.405 36.995 180.865 ;
        RECT 37.205 180.765 37.465 181.155 ;
        RECT 37.655 181.975 38.620 181.985 ;
        RECT 38.790 182.065 38.960 182.445 ;
        RECT 39.550 182.405 39.720 182.695 ;
        RECT 39.900 182.575 40.230 182.955 ;
        RECT 39.550 182.235 40.350 182.405 ;
        RECT 37.655 181.815 38.330 181.975 ;
        RECT 38.790 181.895 40.010 182.065 ;
        RECT 37.655 181.025 37.865 181.815 ;
        RECT 38.790 181.805 38.960 181.895 ;
        RECT 38.035 181.025 38.385 181.645 ;
        RECT 38.555 181.635 38.960 181.805 ;
        RECT 38.555 180.855 38.725 181.635 ;
        RECT 38.895 181.185 39.115 181.465 ;
        RECT 39.295 181.355 39.835 181.725 ;
        RECT 40.180 181.645 40.350 182.235 ;
        RECT 40.570 181.815 40.875 182.955 ;
        RECT 41.045 181.765 41.300 182.645 ;
        RECT 40.180 181.615 40.920 181.645 ;
        RECT 38.895 181.015 39.425 181.185 ;
        RECT 37.205 180.595 37.555 180.765 ;
        RECT 37.775 180.575 38.725 180.855 ;
        RECT 38.895 180.405 39.085 180.845 ;
        RECT 39.255 180.785 39.425 181.015 ;
        RECT 39.595 180.955 39.835 181.355 ;
        RECT 40.005 181.315 40.920 181.615 ;
        RECT 40.005 181.140 40.330 181.315 ;
        RECT 40.005 180.785 40.325 181.140 ;
        RECT 41.090 181.115 41.300 181.765 ;
        RECT 41.935 181.865 43.145 182.955 ;
        RECT 41.935 181.325 42.455 181.865 ;
        RECT 42.625 181.155 43.145 181.695 ;
        RECT 39.255 180.615 40.325 180.785 ;
        RECT 40.570 180.405 40.875 180.865 ;
        RECT 41.045 180.585 41.300 181.115 ;
        RECT 41.935 180.405 43.145 181.155 ;
        RECT 8.270 180.235 43.230 180.405 ;
        RECT 8.355 179.485 9.565 180.235 ;
        RECT 10.255 179.755 10.535 180.235 ;
        RECT 10.705 179.585 10.965 179.975 ;
        RECT 11.140 179.755 11.395 180.235 ;
        RECT 11.565 179.585 11.860 179.975 ;
        RECT 12.040 179.755 12.315 180.235 ;
        RECT 12.485 179.735 12.785 180.065 ;
        RECT 8.355 178.945 8.875 179.485 ;
        RECT 10.210 179.415 11.860 179.585 ;
        RECT 9.045 178.775 9.565 179.315 ;
        RECT 8.355 177.685 9.565 178.775 ;
        RECT 10.210 178.905 10.615 179.415 ;
        RECT 10.785 179.075 11.925 179.245 ;
        RECT 10.210 178.735 10.965 178.905 ;
        RECT 10.250 177.685 10.535 178.555 ;
        RECT 10.705 178.485 10.965 178.735 ;
        RECT 11.755 178.825 11.925 179.075 ;
        RECT 12.095 178.995 12.445 179.565 ;
        RECT 12.615 178.825 12.785 179.735 ;
        RECT 12.975 179.505 13.265 180.235 ;
        RECT 12.965 178.995 13.265 179.325 ;
        RECT 13.445 179.305 13.675 179.945 ;
        RECT 13.855 179.685 14.165 180.055 ;
        RECT 14.345 179.865 15.015 180.235 ;
        RECT 13.855 179.485 15.085 179.685 ;
        RECT 13.445 178.995 13.970 179.305 ;
        RECT 14.150 178.995 14.615 179.305 ;
        RECT 11.755 178.655 12.785 178.825 ;
        RECT 14.795 178.815 15.085 179.485 ;
        RECT 10.705 178.315 11.825 178.485 ;
        RECT 10.705 177.855 10.965 178.315 ;
        RECT 11.140 177.685 11.395 178.145 ;
        RECT 11.565 177.855 11.825 178.315 ;
        RECT 11.995 177.685 12.305 178.485 ;
        RECT 12.475 177.855 12.785 178.655 ;
        RECT 12.975 178.575 14.135 178.815 ;
        RECT 12.975 177.865 13.235 178.575 ;
        RECT 13.405 177.685 13.735 178.395 ;
        RECT 13.905 177.865 14.135 178.575 ;
        RECT 14.315 178.595 15.085 178.815 ;
        RECT 14.315 177.865 14.585 178.595 ;
        RECT 14.765 177.685 15.105 178.415 ;
        RECT 15.275 177.865 15.535 180.055 ;
        RECT 15.805 179.755 16.105 180.235 ;
        RECT 16.275 179.585 16.535 180.040 ;
        RECT 16.705 179.755 16.965 180.235 ;
        RECT 17.145 179.585 17.405 180.040 ;
        RECT 17.575 179.755 17.825 180.235 ;
        RECT 18.005 179.585 18.265 180.040 ;
        RECT 18.435 179.755 18.685 180.235 ;
        RECT 18.865 179.585 19.125 180.040 ;
        RECT 19.295 179.755 19.540 180.235 ;
        RECT 19.710 179.585 19.985 180.040 ;
        RECT 20.155 179.755 20.400 180.235 ;
        RECT 20.570 179.585 20.830 180.040 ;
        RECT 21.000 179.755 21.260 180.235 ;
        RECT 21.430 179.585 21.690 180.040 ;
        RECT 21.860 179.755 22.120 180.235 ;
        RECT 22.290 179.585 22.550 180.040 ;
        RECT 22.720 179.675 22.980 180.235 ;
        RECT 15.805 179.415 22.550 179.585 ;
        RECT 15.805 178.875 16.970 179.415 ;
        RECT 23.150 179.245 23.400 180.055 ;
        RECT 23.580 179.710 23.840 180.235 ;
        RECT 24.010 179.245 24.260 180.055 ;
        RECT 24.440 179.725 24.745 180.235 ;
        RECT 17.140 178.995 24.260 179.245 ;
        RECT 24.430 178.995 24.745 179.555 ;
        RECT 24.920 179.495 25.175 180.065 ;
        RECT 25.345 179.835 25.675 180.235 ;
        RECT 26.100 179.700 26.630 180.065 ;
        RECT 26.820 179.895 27.095 180.065 ;
        RECT 26.815 179.725 27.095 179.895 ;
        RECT 26.100 179.665 26.275 179.700 ;
        RECT 25.345 179.495 26.275 179.665 ;
        RECT 15.775 178.825 16.970 178.875 ;
        RECT 15.775 178.705 22.550 178.825 ;
        RECT 15.805 178.600 22.550 178.705 ;
        RECT 15.805 177.685 16.075 178.430 ;
        RECT 16.245 177.860 16.535 178.600 ;
        RECT 17.145 178.585 22.550 178.600 ;
        RECT 16.705 177.690 16.960 178.415 ;
        RECT 17.145 177.860 17.405 178.585 ;
        RECT 17.575 177.690 17.820 178.415 ;
        RECT 18.005 177.860 18.265 178.585 ;
        RECT 18.435 177.690 18.680 178.415 ;
        RECT 18.865 177.860 19.125 178.585 ;
        RECT 19.295 177.690 19.540 178.415 ;
        RECT 19.710 177.860 19.970 178.585 ;
        RECT 20.140 177.690 20.400 178.415 ;
        RECT 20.570 177.860 20.830 178.585 ;
        RECT 21.000 177.690 21.260 178.415 ;
        RECT 21.430 177.860 21.690 178.585 ;
        RECT 21.860 177.690 22.120 178.415 ;
        RECT 22.290 177.860 22.550 178.585 ;
        RECT 22.720 177.690 22.980 178.485 ;
        RECT 23.150 177.860 23.400 178.995 ;
        RECT 16.705 177.685 22.980 177.690 ;
        RECT 23.580 177.685 23.840 178.495 ;
        RECT 24.015 177.855 24.260 178.995 ;
        RECT 24.920 178.825 25.090 179.495 ;
        RECT 25.345 179.325 25.515 179.495 ;
        RECT 25.260 178.995 25.515 179.325 ;
        RECT 25.740 178.995 25.935 179.325 ;
        RECT 24.440 177.685 24.735 178.495 ;
        RECT 24.920 177.855 25.255 178.825 ;
        RECT 25.425 177.685 25.595 178.825 ;
        RECT 25.765 178.025 25.935 178.995 ;
        RECT 26.105 178.365 26.275 179.495 ;
        RECT 26.445 178.705 26.615 179.505 ;
        RECT 26.820 178.905 27.095 179.725 ;
        RECT 27.265 178.705 27.455 180.065 ;
        RECT 27.635 179.700 28.145 180.235 ;
        RECT 28.365 179.425 28.610 180.030 ;
        RECT 29.170 179.605 29.455 180.065 ;
        RECT 29.625 179.775 29.895 180.235 ;
        RECT 29.170 179.435 30.125 179.605 ;
        RECT 27.655 179.255 28.885 179.425 ;
        RECT 26.445 178.535 27.455 178.705 ;
        RECT 27.625 178.690 28.375 178.880 ;
        RECT 26.105 178.195 27.230 178.365 ;
        RECT 27.625 178.025 27.795 178.690 ;
        RECT 28.545 178.445 28.885 179.255 ;
        RECT 29.055 178.705 29.745 179.265 ;
        RECT 29.915 178.535 30.125 179.435 ;
        RECT 25.765 177.855 27.795 178.025 ;
        RECT 27.965 177.685 28.135 178.445 ;
        RECT 28.370 178.035 28.885 178.445 ;
        RECT 29.170 178.315 30.125 178.535 ;
        RECT 30.295 179.265 30.695 180.065 ;
        RECT 30.885 179.605 31.165 180.065 ;
        RECT 31.685 179.775 32.010 180.235 ;
        RECT 30.885 179.435 32.010 179.605 ;
        RECT 32.180 179.495 32.565 180.065 ;
        RECT 31.560 179.325 32.010 179.435 ;
        RECT 30.295 178.705 31.390 179.265 ;
        RECT 31.560 178.995 32.115 179.325 ;
        RECT 29.170 177.855 29.455 178.315 ;
        RECT 29.625 177.685 29.895 178.145 ;
        RECT 30.295 177.855 30.695 178.705 ;
        RECT 31.560 178.535 32.010 178.995 ;
        RECT 32.285 178.825 32.565 179.495 ;
        RECT 32.735 179.485 33.945 180.235 ;
        RECT 34.115 179.510 34.405 180.235 ;
        RECT 32.735 178.945 33.255 179.485 ;
        RECT 30.885 178.315 32.010 178.535 ;
        RECT 30.885 177.855 31.165 178.315 ;
        RECT 31.685 177.685 32.010 178.145 ;
        RECT 32.180 177.855 32.565 178.825 ;
        RECT 33.425 178.775 33.945 179.315 ;
        RECT 35.495 179.290 35.835 180.065 ;
        RECT 36.005 179.775 36.175 180.235 ;
        RECT 36.415 179.800 36.775 180.065 ;
        RECT 36.415 179.795 36.770 179.800 ;
        RECT 36.415 179.785 36.765 179.795 ;
        RECT 36.415 179.780 36.760 179.785 ;
        RECT 36.415 179.770 36.755 179.780 ;
        RECT 37.405 179.775 37.575 180.235 ;
        RECT 36.415 179.765 36.750 179.770 ;
        RECT 36.415 179.755 36.740 179.765 ;
        RECT 36.415 179.745 36.730 179.755 ;
        RECT 36.415 179.605 36.715 179.745 ;
        RECT 36.005 179.415 36.715 179.605 ;
        RECT 36.905 179.605 37.235 179.685 ;
        RECT 37.745 179.605 38.085 180.065 ;
        RECT 36.905 179.415 38.085 179.605 ;
        RECT 38.255 179.735 38.515 180.065 ;
        RECT 38.685 179.875 39.015 180.235 ;
        RECT 39.270 179.855 40.570 180.065 ;
        RECT 38.255 179.725 38.485 179.735 ;
        RECT 32.735 177.685 33.945 178.775 ;
        RECT 34.115 177.685 34.405 178.850 ;
        RECT 35.495 177.855 35.775 179.290 ;
        RECT 36.005 178.845 36.290 179.415 ;
        RECT 36.475 179.015 36.945 179.245 ;
        RECT 37.115 179.225 37.445 179.245 ;
        RECT 37.115 179.045 37.565 179.225 ;
        RECT 37.755 179.045 38.085 179.245 ;
        RECT 36.005 178.630 37.155 178.845 ;
        RECT 35.945 177.685 36.655 178.460 ;
        RECT 36.825 177.855 37.155 178.630 ;
        RECT 37.350 177.930 37.565 179.045 ;
        RECT 37.855 178.705 38.085 179.045 ;
        RECT 38.255 178.535 38.425 179.725 ;
        RECT 39.270 179.705 39.440 179.855 ;
        RECT 38.685 179.580 39.440 179.705 ;
        RECT 38.595 179.535 39.440 179.580 ;
        RECT 38.595 179.415 38.865 179.535 ;
        RECT 38.595 178.840 38.765 179.415 ;
        RECT 38.995 178.975 39.405 179.280 ;
        RECT 39.695 179.245 39.905 179.645 ;
        RECT 39.575 179.035 39.905 179.245 ;
        RECT 40.150 179.245 40.370 179.645 ;
        RECT 40.845 179.470 41.300 180.235 ;
        RECT 41.935 179.485 43.145 180.235 ;
        RECT 40.150 179.035 40.625 179.245 ;
        RECT 40.815 179.045 41.305 179.245 ;
        RECT 38.595 178.805 38.795 178.840 ;
        RECT 40.125 178.805 41.300 178.865 ;
        RECT 38.595 178.695 41.300 178.805 ;
        RECT 38.655 178.635 40.455 178.695 ;
        RECT 40.125 178.605 40.455 178.635 ;
        RECT 37.745 177.685 38.075 178.405 ;
        RECT 38.255 177.855 38.515 178.535 ;
        RECT 38.685 177.685 38.935 178.465 ;
        RECT 39.185 178.435 40.020 178.445 ;
        RECT 40.610 178.435 40.795 178.525 ;
        RECT 39.185 178.235 40.795 178.435 ;
        RECT 39.185 177.855 39.435 178.235 ;
        RECT 40.565 178.195 40.795 178.235 ;
        RECT 41.045 178.075 41.300 178.695 ;
        RECT 39.605 177.685 39.960 178.065 ;
        RECT 40.965 177.855 41.300 178.075 ;
        RECT 41.935 178.775 42.455 179.315 ;
        RECT 42.625 178.945 43.145 179.485 ;
        RECT 41.935 177.685 43.145 178.775 ;
        RECT 8.270 177.515 43.230 177.685 ;
        RECT 8.355 176.425 9.565 177.515 ;
        RECT 9.735 176.425 11.405 177.515 ;
        RECT 12.040 176.845 12.295 177.345 ;
        RECT 12.465 177.015 12.795 177.515 ;
        RECT 12.040 176.675 12.790 176.845 ;
        RECT 8.355 175.715 8.875 176.255 ;
        RECT 9.045 175.885 9.565 176.425 ;
        RECT 9.735 175.735 10.485 176.255 ;
        RECT 10.655 175.905 11.405 176.425 ;
        RECT 12.040 175.855 12.390 176.505 ;
        RECT 8.355 174.965 9.565 175.715 ;
        RECT 9.735 174.965 11.405 175.735 ;
        RECT 12.560 175.685 12.790 176.675 ;
        RECT 12.040 175.515 12.790 175.685 ;
        RECT 12.040 175.225 12.295 175.515 ;
        RECT 12.465 174.965 12.795 175.345 ;
        RECT 12.965 175.225 13.135 177.345 ;
        RECT 13.305 176.545 13.630 177.330 ;
        RECT 13.800 177.055 14.050 177.515 ;
        RECT 14.220 177.015 14.470 177.345 ;
        RECT 14.685 177.015 15.365 177.345 ;
        RECT 14.220 176.885 14.390 177.015 ;
        RECT 13.995 176.715 14.390 176.885 ;
        RECT 13.365 175.495 13.825 176.545 ;
        RECT 13.995 175.355 14.165 176.715 ;
        RECT 14.560 176.455 15.025 176.845 ;
        RECT 14.335 175.645 14.685 176.265 ;
        RECT 14.855 175.865 15.025 176.455 ;
        RECT 15.195 176.235 15.365 177.015 ;
        RECT 15.535 176.915 15.705 177.255 ;
        RECT 15.940 177.085 16.270 177.515 ;
        RECT 16.440 176.915 16.610 177.255 ;
        RECT 16.905 177.055 17.275 177.515 ;
        RECT 15.535 176.745 16.610 176.915 ;
        RECT 17.445 176.885 17.615 177.345 ;
        RECT 17.850 177.005 18.720 177.345 ;
        RECT 18.890 177.055 19.140 177.515 ;
        RECT 17.055 176.715 17.615 176.885 ;
        RECT 17.055 176.575 17.225 176.715 ;
        RECT 15.725 176.405 17.225 176.575 ;
        RECT 17.920 176.545 18.380 176.835 ;
        RECT 15.195 176.065 16.885 176.235 ;
        RECT 14.855 175.645 15.210 175.865 ;
        RECT 15.380 175.355 15.550 176.065 ;
        RECT 15.755 175.645 16.545 175.895 ;
        RECT 16.715 175.885 16.885 176.065 ;
        RECT 17.055 175.715 17.225 176.405 ;
        RECT 13.495 174.965 13.825 175.325 ;
        RECT 13.995 175.185 14.490 175.355 ;
        RECT 14.695 175.185 15.550 175.355 ;
        RECT 16.425 174.965 16.755 175.425 ;
        RECT 16.965 175.325 17.225 175.715 ;
        RECT 17.415 176.535 18.380 176.545 ;
        RECT 18.550 176.625 18.720 177.005 ;
        RECT 19.310 176.965 19.480 177.255 ;
        RECT 19.660 177.135 19.990 177.515 ;
        RECT 19.310 176.795 20.110 176.965 ;
        RECT 17.415 176.375 18.090 176.535 ;
        RECT 18.550 176.455 19.770 176.625 ;
        RECT 17.415 175.585 17.625 176.375 ;
        RECT 18.550 176.365 18.720 176.455 ;
        RECT 17.795 175.585 18.145 176.205 ;
        RECT 18.315 176.195 18.720 176.365 ;
        RECT 18.315 175.415 18.485 176.195 ;
        RECT 18.655 175.745 18.875 176.025 ;
        RECT 19.055 175.915 19.595 176.285 ;
        RECT 19.940 176.205 20.110 176.795 ;
        RECT 20.330 176.375 20.635 177.515 ;
        RECT 20.805 176.325 21.060 177.205 ;
        RECT 21.235 176.350 21.525 177.515 ;
        RECT 21.695 176.795 22.155 177.345 ;
        RECT 22.345 176.795 22.675 177.515 ;
        RECT 19.940 176.175 20.680 176.205 ;
        RECT 18.655 175.575 19.185 175.745 ;
        RECT 16.965 175.155 17.315 175.325 ;
        RECT 17.535 175.135 18.485 175.415 ;
        RECT 18.655 174.965 18.845 175.405 ;
        RECT 19.015 175.345 19.185 175.575 ;
        RECT 19.355 175.515 19.595 175.915 ;
        RECT 19.765 175.875 20.680 176.175 ;
        RECT 19.765 175.700 20.090 175.875 ;
        RECT 19.765 175.345 20.085 175.700 ;
        RECT 20.850 175.675 21.060 176.325 ;
        RECT 19.015 175.175 20.085 175.345 ;
        RECT 20.330 174.965 20.635 175.425 ;
        RECT 20.805 175.145 21.060 175.675 ;
        RECT 21.235 174.965 21.525 175.690 ;
        RECT 21.695 175.425 21.945 176.795 ;
        RECT 22.875 176.625 23.175 177.175 ;
        RECT 23.345 176.845 23.625 177.515 ;
        RECT 22.235 176.455 23.175 176.625 ;
        RECT 22.235 176.205 22.405 176.455 ;
        RECT 23.545 176.205 23.810 176.565 ;
        RECT 22.115 175.875 22.405 176.205 ;
        RECT 22.575 175.955 22.915 176.205 ;
        RECT 23.135 175.955 23.810 176.205 ;
        RECT 23.995 176.545 24.305 177.345 ;
        RECT 24.475 176.715 24.785 177.515 ;
        RECT 24.955 176.885 25.215 177.345 ;
        RECT 25.385 177.055 25.640 177.515 ;
        RECT 25.815 176.885 26.075 177.345 ;
        RECT 24.955 176.715 26.075 176.885 ;
        RECT 23.995 176.375 25.025 176.545 ;
        RECT 22.235 175.785 22.405 175.875 ;
        RECT 22.235 175.595 23.625 175.785 ;
        RECT 21.695 175.135 22.255 175.425 ;
        RECT 22.425 174.965 22.675 175.425 ;
        RECT 23.295 175.235 23.625 175.595 ;
        RECT 23.995 175.465 24.165 176.375 ;
        RECT 24.335 175.635 24.685 176.205 ;
        RECT 24.855 176.125 25.025 176.375 ;
        RECT 25.815 176.465 26.075 176.715 ;
        RECT 26.245 176.645 26.530 177.515 ;
        RECT 26.810 176.645 27.095 177.515 ;
        RECT 27.265 176.885 27.525 177.345 ;
        RECT 27.700 177.055 27.955 177.515 ;
        RECT 28.125 176.885 28.385 177.345 ;
        RECT 27.265 176.715 28.385 176.885 ;
        RECT 28.555 176.715 28.865 177.515 ;
        RECT 27.265 176.465 27.525 176.715 ;
        RECT 29.035 176.545 29.345 177.345 ;
        RECT 25.815 176.295 26.570 176.465 ;
        RECT 24.855 175.955 25.995 176.125 ;
        RECT 26.165 175.785 26.570 176.295 ;
        RECT 24.920 175.615 26.570 175.785 ;
        RECT 26.770 176.295 27.525 176.465 ;
        RECT 28.315 176.375 29.345 176.545 ;
        RECT 26.770 175.785 27.175 176.295 ;
        RECT 28.315 176.125 28.485 176.375 ;
        RECT 27.345 175.955 28.485 176.125 ;
        RECT 26.770 175.615 28.420 175.785 ;
        RECT 28.655 175.635 29.005 176.205 ;
        RECT 23.995 175.135 24.295 175.465 ;
        RECT 24.465 174.965 24.740 175.445 ;
        RECT 24.920 175.225 25.215 175.615 ;
        RECT 25.385 174.965 25.640 175.445 ;
        RECT 25.815 175.225 26.075 175.615 ;
        RECT 26.245 174.965 26.525 175.445 ;
        RECT 26.815 174.965 27.095 175.445 ;
        RECT 27.265 175.225 27.525 175.615 ;
        RECT 27.700 174.965 27.955 175.445 ;
        RECT 28.125 175.225 28.420 175.615 ;
        RECT 29.175 175.465 29.345 176.375 ;
        RECT 28.600 174.965 28.875 175.445 ;
        RECT 29.045 175.135 29.345 175.465 ;
        RECT 29.515 175.910 29.795 177.345 ;
        RECT 29.965 176.740 30.675 177.515 ;
        RECT 30.845 176.570 31.175 177.345 ;
        RECT 30.025 176.355 31.175 176.570 ;
        RECT 29.515 175.135 29.855 175.910 ;
        RECT 30.025 175.785 30.310 176.355 ;
        RECT 30.495 175.955 30.965 176.185 ;
        RECT 31.370 176.155 31.585 177.270 ;
        RECT 31.765 176.795 32.095 177.515 ;
        RECT 31.875 176.155 32.105 176.495 ;
        RECT 32.275 176.425 33.945 177.515 ;
        RECT 31.135 175.975 31.585 176.155 ;
        RECT 31.135 175.955 31.465 175.975 ;
        RECT 31.775 175.955 32.105 176.155 ;
        RECT 30.025 175.595 30.735 175.785 ;
        RECT 30.435 175.455 30.735 175.595 ;
        RECT 30.925 175.595 32.105 175.785 ;
        RECT 30.925 175.515 31.255 175.595 ;
        RECT 30.435 175.445 30.750 175.455 ;
        RECT 30.435 175.435 30.760 175.445 ;
        RECT 30.435 175.430 30.770 175.435 ;
        RECT 30.025 174.965 30.195 175.425 ;
        RECT 30.435 175.420 30.775 175.430 ;
        RECT 30.435 175.415 30.780 175.420 ;
        RECT 30.435 175.405 30.785 175.415 ;
        RECT 30.435 175.400 30.790 175.405 ;
        RECT 30.435 175.135 30.795 175.400 ;
        RECT 31.425 174.965 31.595 175.425 ;
        RECT 31.765 175.135 32.105 175.595 ;
        RECT 32.275 175.735 33.025 176.255 ;
        RECT 33.195 175.905 33.945 176.425 ;
        RECT 34.115 176.350 34.405 177.515 ;
        RECT 34.575 176.545 34.885 177.345 ;
        RECT 35.055 176.715 35.365 177.515 ;
        RECT 35.535 176.885 35.795 177.345 ;
        RECT 35.965 177.055 36.220 177.515 ;
        RECT 36.395 176.885 36.655 177.345 ;
        RECT 35.535 176.715 36.655 176.885 ;
        RECT 34.575 176.375 35.605 176.545 ;
        RECT 32.275 174.965 33.945 175.735 ;
        RECT 34.115 174.965 34.405 175.690 ;
        RECT 34.575 175.465 34.745 176.375 ;
        RECT 34.915 175.635 35.265 176.205 ;
        RECT 35.435 176.125 35.605 176.375 ;
        RECT 36.395 176.465 36.655 176.715 ;
        RECT 36.825 176.645 37.110 177.515 ;
        RECT 37.335 176.545 37.645 177.345 ;
        RECT 37.815 176.715 38.125 177.515 ;
        RECT 38.295 176.885 38.555 177.345 ;
        RECT 38.725 177.055 38.980 177.515 ;
        RECT 39.155 176.885 39.415 177.345 ;
        RECT 38.295 176.715 39.415 176.885 ;
        RECT 36.395 176.295 37.150 176.465 ;
        RECT 35.435 175.955 36.575 176.125 ;
        RECT 36.745 175.785 37.150 176.295 ;
        RECT 35.500 175.615 37.150 175.785 ;
        RECT 37.335 176.375 38.365 176.545 ;
        RECT 34.575 175.135 34.875 175.465 ;
        RECT 35.045 174.965 35.320 175.445 ;
        RECT 35.500 175.225 35.795 175.615 ;
        RECT 35.965 174.965 36.220 175.445 ;
        RECT 36.395 175.225 36.655 175.615 ;
        RECT 37.335 175.465 37.505 176.375 ;
        RECT 37.675 175.635 38.025 176.205 ;
        RECT 38.195 176.125 38.365 176.375 ;
        RECT 39.155 176.465 39.415 176.715 ;
        RECT 39.585 176.645 39.870 177.515 ;
        RECT 39.155 176.295 39.910 176.465 ;
        RECT 40.095 176.425 41.765 177.515 ;
        RECT 38.195 175.955 39.335 176.125 ;
        RECT 39.505 175.785 39.910 176.295 ;
        RECT 38.260 175.615 39.910 175.785 ;
        RECT 40.095 175.735 40.845 176.255 ;
        RECT 41.015 175.905 41.765 176.425 ;
        RECT 41.935 176.425 43.145 177.515 ;
        RECT 41.935 175.885 42.455 176.425 ;
        RECT 36.825 174.965 37.105 175.445 ;
        RECT 37.335 175.135 37.635 175.465 ;
        RECT 37.805 174.965 38.080 175.445 ;
        RECT 38.260 175.225 38.555 175.615 ;
        RECT 38.725 174.965 38.980 175.445 ;
        RECT 39.155 175.225 39.415 175.615 ;
        RECT 39.585 174.965 39.865 175.445 ;
        RECT 40.095 174.965 41.765 175.735 ;
        RECT 42.625 175.715 43.145 176.255 ;
        RECT 41.935 174.965 43.145 175.715 ;
        RECT 8.270 174.795 43.230 174.965 ;
        RECT 58.955 160.995 60.905 161.165 ;
        RECT 58.955 158.660 59.125 160.995 ;
        RECT 59.755 160.485 60.105 160.655 ;
        RECT 57.305 158.490 59.130 158.660 ;
        RECT 57.645 157.350 57.855 158.490 ;
        RECT 58.525 158.485 59.130 158.490 ;
        RECT 58.025 157.400 58.355 158.320 ;
        RECT 58.955 157.505 59.125 158.485 ;
        RECT 59.525 158.230 59.695 160.270 ;
        RECT 60.165 158.230 60.335 160.270 ;
        RECT 59.755 157.845 60.105 158.015 ;
        RECT 60.735 157.505 60.905 160.995 ;
        RECT 58.025 157.340 58.770 157.400 ;
        RECT 58.125 157.230 58.770 157.340 ;
        RECT 58.955 157.335 60.905 157.505 ;
        RECT 57.625 157.115 57.955 157.170 ;
        RECT 57.165 156.935 57.955 157.115 ;
        RECT 57.625 156.930 57.955 156.935 ;
        RECT 57.625 155.940 57.855 156.760 ;
        RECT 58.125 156.740 58.355 157.230 ;
        RECT 58.025 156.110 58.355 156.740 ;
        RECT 59.065 156.735 60.815 156.905 ;
        RECT 59.065 155.955 59.235 156.735 ;
        RECT 59.775 156.225 60.105 156.395 ;
        RECT 58.525 155.940 59.240 155.955 ;
        RECT 57.305 155.780 59.240 155.940 ;
        RECT 57.305 155.770 58.685 155.780 ;
        RECT 59.065 154.915 59.235 155.780 ;
        RECT 59.635 155.595 59.805 156.055 ;
        RECT 60.075 155.595 60.245 156.055 ;
        RECT 59.775 155.255 60.105 155.425 ;
        RECT 60.645 154.915 60.815 156.735 ;
        RECT 59.065 154.745 60.815 154.915 ;
        RECT 58.790 131.165 60.740 131.335 ;
        RECT 58.790 128.830 58.960 131.165 ;
        RECT 59.590 130.655 59.940 130.825 ;
        RECT 57.140 128.660 58.965 128.830 ;
        RECT 57.480 127.520 57.690 128.660 ;
        RECT 58.360 128.655 58.965 128.660 ;
        RECT 57.860 127.570 58.190 128.490 ;
        RECT 58.790 127.675 58.960 128.655 ;
        RECT 59.360 128.400 59.530 130.440 ;
        RECT 60.000 128.400 60.170 130.440 ;
        RECT 59.590 128.015 59.940 128.185 ;
        RECT 60.570 127.675 60.740 131.165 ;
        RECT 57.860 127.510 58.605 127.570 ;
        RECT 57.960 127.400 58.605 127.510 ;
        RECT 58.790 127.505 60.740 127.675 ;
        RECT 57.460 127.285 57.790 127.340 ;
        RECT 57.000 127.105 57.790 127.285 ;
        RECT 57.460 127.100 57.790 127.105 ;
        RECT 57.460 126.110 57.690 126.930 ;
        RECT 57.960 126.910 58.190 127.400 ;
        RECT 57.860 126.280 58.190 126.910 ;
        RECT 58.900 126.905 60.650 127.075 ;
        RECT 58.900 126.125 59.070 126.905 ;
        RECT 59.610 126.395 59.940 126.565 ;
        RECT 58.360 126.110 59.075 126.125 ;
        RECT 57.140 125.950 59.075 126.110 ;
        RECT 57.140 125.940 58.520 125.950 ;
        RECT 58.900 125.085 59.070 125.950 ;
        RECT 59.470 125.765 59.640 126.225 ;
        RECT 59.910 125.765 60.080 126.225 ;
        RECT 59.610 125.425 59.940 125.595 ;
        RECT 60.480 125.085 60.650 126.905 ;
        RECT 58.900 124.915 60.650 125.085 ;
        RECT 19.900 104.560 21.850 104.730 ;
        RECT 19.900 102.225 20.070 104.560 ;
        RECT 20.700 104.050 21.050 104.220 ;
        RECT 18.250 102.055 20.075 102.225 ;
        RECT 18.590 100.915 18.800 102.055 ;
        RECT 19.470 102.050 20.075 102.055 ;
        RECT 18.970 100.965 19.300 101.885 ;
        RECT 19.900 101.070 20.070 102.050 ;
        RECT 20.470 101.795 20.640 103.835 ;
        RECT 21.110 101.795 21.280 103.835 ;
        RECT 20.700 101.410 21.050 101.580 ;
        RECT 21.680 101.070 21.850 104.560 ;
        RECT 34.960 102.900 37.120 103.070 ;
        RECT 34.960 101.525 35.130 102.900 ;
        RECT 35.470 102.030 35.640 102.360 ;
        RECT 35.810 102.330 36.270 102.500 ;
        RECT 35.810 101.890 36.270 102.060 ;
        RECT 36.440 102.030 36.610 102.360 ;
        RECT 33.835 101.490 35.165 101.525 ;
        RECT 36.950 101.490 37.120 102.900 ;
        RECT 33.835 101.470 37.120 101.490 ;
        RECT 40.000 102.890 42.160 103.060 ;
        RECT 40.000 101.480 40.170 102.890 ;
        RECT 40.510 102.020 40.680 102.350 ;
        RECT 40.850 102.320 41.310 102.490 ;
        RECT 40.850 101.880 41.310 102.050 ;
        RECT 41.480 102.020 41.650 102.350 ;
        RECT 41.990 101.480 42.160 102.890 ;
        RECT 40.000 101.470 42.160 101.480 ;
        RECT 44.960 102.880 47.120 103.050 ;
        RECT 44.960 101.470 45.130 102.880 ;
        RECT 45.470 102.010 45.640 102.340 ;
        RECT 45.810 102.310 46.270 102.480 ;
        RECT 45.810 101.870 46.270 102.040 ;
        RECT 46.440 102.010 46.610 102.340 ;
        RECT 46.950 101.470 47.120 102.880 ;
        RECT 33.835 101.300 47.120 101.470 ;
        RECT 33.835 101.285 35.165 101.300 ;
        RECT 18.970 100.905 19.715 100.965 ;
        RECT 19.070 100.795 19.715 100.905 ;
        RECT 19.900 100.900 21.850 101.070 ;
        RECT 38.585 100.955 38.755 101.300 ;
        RECT 43.340 100.920 43.510 101.300 ;
        RECT 18.570 100.680 18.900 100.735 ;
        RECT 18.110 100.500 18.900 100.680 ;
        RECT 18.570 100.495 18.900 100.500 ;
        RECT 18.570 99.505 18.800 100.325 ;
        RECT 19.070 100.305 19.300 100.795 ;
        RECT 18.970 99.675 19.300 100.305 ;
        RECT 20.010 100.300 21.760 100.470 ;
        RECT 20.010 99.520 20.180 100.300 ;
        RECT 20.720 99.790 21.050 99.960 ;
        RECT 19.470 99.505 20.185 99.520 ;
        RECT 18.250 99.345 20.185 99.505 ;
        RECT 18.250 99.335 19.630 99.345 ;
        RECT 20.010 98.480 20.180 99.345 ;
        RECT 20.580 99.160 20.750 99.620 ;
        RECT 21.020 99.160 21.190 99.620 ;
        RECT 20.720 98.820 21.050 98.990 ;
        RECT 21.590 98.480 21.760 100.300 ;
        RECT 20.010 98.310 21.760 98.480 ;
        RECT 21.590 97.670 21.760 98.310 ;
        RECT 59.250 100.305 61.200 100.475 ;
        RECT 59.250 97.970 59.420 100.305 ;
        RECT 60.050 99.795 60.400 99.965 ;
        RECT 57.600 97.800 59.425 97.970 ;
        RECT 57.940 96.660 58.150 97.800 ;
        RECT 58.820 97.795 59.425 97.800 ;
        RECT 58.320 96.710 58.650 97.630 ;
        RECT 59.250 96.815 59.420 97.795 ;
        RECT 59.820 97.540 59.990 99.580 ;
        RECT 60.460 97.540 60.630 99.580 ;
        RECT 60.050 97.155 60.400 97.325 ;
        RECT 61.030 96.815 61.200 100.305 ;
        RECT 58.320 96.650 59.065 96.710 ;
        RECT 58.420 96.540 59.065 96.650 ;
        RECT 59.250 96.645 61.200 96.815 ;
        RECT 57.920 96.425 58.250 96.480 ;
        RECT 57.460 96.245 58.250 96.425 ;
        RECT 57.920 96.240 58.250 96.245 ;
        RECT 57.920 95.250 58.150 96.070 ;
        RECT 58.420 96.050 58.650 96.540 ;
        RECT 58.320 95.420 58.650 96.050 ;
        RECT 59.360 96.045 61.110 96.215 ;
        RECT 59.360 95.265 59.530 96.045 ;
        RECT 60.070 95.535 60.400 95.705 ;
        RECT 58.820 95.250 59.535 95.265 ;
        RECT 57.600 95.090 59.535 95.250 ;
        RECT 57.600 95.080 58.980 95.090 ;
        RECT 59.360 94.225 59.530 95.090 ;
        RECT 59.930 94.905 60.100 95.365 ;
        RECT 60.370 94.905 60.540 95.365 ;
        RECT 60.070 94.565 60.400 94.735 ;
        RECT 60.940 94.225 61.110 96.045 ;
        RECT 59.360 94.055 61.110 94.225 ;
        RECT 20.050 93.490 22.000 93.660 ;
        RECT 20.050 91.155 20.220 93.490 ;
        RECT 20.850 92.980 21.200 93.150 ;
        RECT 18.400 90.985 20.225 91.155 ;
        RECT 18.740 89.845 18.950 90.985 ;
        RECT 19.620 90.980 20.225 90.985 ;
        RECT 19.120 89.895 19.450 90.815 ;
        RECT 20.050 90.000 20.220 90.980 ;
        RECT 20.620 90.725 20.790 92.765 ;
        RECT 21.260 90.725 21.430 92.765 ;
        RECT 20.850 90.340 21.200 90.510 ;
        RECT 21.830 90.000 22.000 93.490 ;
        RECT 19.120 89.835 19.865 89.895 ;
        RECT 19.220 89.725 19.865 89.835 ;
        RECT 20.050 89.830 22.000 90.000 ;
        RECT 18.720 89.610 19.050 89.665 ;
        RECT 18.260 89.430 19.050 89.610 ;
        RECT 18.720 89.425 19.050 89.430 ;
        RECT 18.720 88.435 18.950 89.255 ;
        RECT 19.220 89.235 19.450 89.725 ;
        RECT 19.120 88.605 19.450 89.235 ;
        RECT 20.160 89.230 21.910 89.400 ;
        RECT 20.160 88.450 20.330 89.230 ;
        RECT 20.870 88.720 21.200 88.890 ;
        RECT 19.620 88.435 20.335 88.450 ;
        RECT 18.400 88.275 20.335 88.435 ;
        RECT 18.400 88.265 19.780 88.275 ;
        RECT 20.160 87.410 20.330 88.275 ;
        RECT 20.730 88.090 20.900 88.550 ;
        RECT 21.170 88.090 21.340 88.550 ;
        RECT 20.870 87.750 21.200 87.920 ;
        RECT 21.740 87.410 21.910 89.230 ;
        RECT 20.160 87.240 21.910 87.410 ;
        RECT 21.725 86.515 21.895 87.240 ;
        RECT 20.000 82.360 21.950 82.530 ;
        RECT 20.000 80.025 20.170 82.360 ;
        RECT 20.800 81.850 21.150 82.020 ;
        RECT 18.350 79.855 20.175 80.025 ;
        RECT 18.690 78.715 18.900 79.855 ;
        RECT 19.570 79.850 20.175 79.855 ;
        RECT 19.070 78.765 19.400 79.685 ;
        RECT 20.000 78.870 20.170 79.850 ;
        RECT 20.570 79.595 20.740 81.635 ;
        RECT 21.210 79.595 21.380 81.635 ;
        RECT 20.800 79.210 21.150 79.380 ;
        RECT 21.780 78.870 21.950 82.360 ;
        RECT 34.755 79.730 34.925 80.055 ;
        RECT 28.765 79.675 36.645 79.730 ;
        RECT 28.765 79.660 39.145 79.675 ;
        RECT 43.310 79.660 46.140 79.675 ;
        RECT 28.765 79.560 46.140 79.660 ;
        RECT 27.040 79.315 28.420 79.325 ;
        RECT 28.765 79.315 28.935 79.560 ;
        RECT 27.040 79.155 28.940 79.315 ;
        RECT 19.070 78.705 19.815 78.765 ;
        RECT 19.170 78.595 19.815 78.705 ;
        RECT 20.000 78.700 21.950 78.870 ;
        RECT 18.670 78.480 19.000 78.535 ;
        RECT 18.210 78.300 19.000 78.480 ;
        RECT 18.670 78.295 19.000 78.300 ;
        RECT 18.670 77.305 18.900 78.125 ;
        RECT 19.170 78.105 19.400 78.595 ;
        RECT 19.070 77.475 19.400 78.105 ;
        RECT 20.110 78.100 21.860 78.270 ;
        RECT 20.110 77.320 20.280 78.100 ;
        RECT 20.820 77.590 21.150 77.760 ;
        RECT 19.570 77.305 20.285 77.320 ;
        RECT 18.350 77.145 20.285 77.305 ;
        RECT 18.350 77.135 19.730 77.145 ;
        RECT 20.110 76.280 20.280 77.145 ;
        RECT 20.680 76.960 20.850 77.420 ;
        RECT 21.120 76.960 21.290 77.420 ;
        RECT 20.820 76.620 21.150 76.790 ;
        RECT 21.690 76.340 21.860 78.100 ;
        RECT 27.380 78.015 27.590 79.155 ;
        RECT 28.260 79.140 28.940 79.155 ;
        RECT 27.760 78.075 28.090 78.985 ;
        RECT 28.765 78.150 28.935 79.140 ;
        RECT 29.275 78.690 29.445 79.020 ;
        RECT 29.660 78.990 30.700 79.160 ;
        RECT 29.660 78.550 30.700 78.720 ;
        RECT 30.915 78.690 31.085 79.020 ;
        RECT 31.425 78.150 31.595 79.560 ;
        RECT 36.315 79.505 46.140 79.560 ;
        RECT 34.590 79.260 35.970 79.270 ;
        RECT 36.315 79.260 36.485 79.505 ;
        RECT 38.830 79.490 43.480 79.505 ;
        RECT 34.590 79.100 36.490 79.260 ;
        RECT 27.760 78.005 28.515 78.075 ;
        RECT 27.860 77.885 28.515 78.005 ;
        RECT 28.765 77.980 31.595 78.150 ;
        RECT 34.930 77.960 35.140 79.100 ;
        RECT 35.810 79.085 36.490 79.100 ;
        RECT 35.310 78.020 35.640 78.930 ;
        RECT 36.315 78.095 36.485 79.085 ;
        RECT 36.825 78.635 36.995 78.965 ;
        RECT 37.210 78.935 38.250 79.105 ;
        RECT 37.210 78.495 38.250 78.665 ;
        RECT 38.465 78.635 38.635 78.965 ;
        RECT 38.975 78.095 39.145 79.490 ;
        RECT 41.585 79.260 42.965 79.270 ;
        RECT 43.310 79.260 43.480 79.490 ;
        RECT 41.585 79.100 43.485 79.260 ;
        RECT 35.310 77.950 36.065 78.020 ;
        RECT 27.360 77.805 27.690 77.835 ;
        RECT 26.990 77.620 27.690 77.805 ;
        RECT 27.360 77.595 27.690 77.620 ;
        RECT 27.360 76.605 27.590 77.425 ;
        RECT 27.860 77.405 28.090 77.885 ;
        RECT 35.410 77.830 36.065 77.950 ;
        RECT 36.315 77.925 39.145 78.095 ;
        RECT 41.925 77.960 42.135 79.100 ;
        RECT 42.805 79.085 43.485 79.100 ;
        RECT 42.305 78.020 42.635 78.930 ;
        RECT 43.310 78.095 43.480 79.085 ;
        RECT 43.820 78.635 43.990 78.965 ;
        RECT 44.205 78.935 45.245 79.105 ;
        RECT 44.205 78.495 45.245 78.665 ;
        RECT 45.460 78.635 45.630 78.965 ;
        RECT 45.970 78.095 46.140 79.505 ;
        RECT 42.305 77.950 43.060 78.020 ;
        RECT 42.405 77.830 43.060 77.950 ;
        RECT 43.310 77.925 46.140 78.095 ;
        RECT 34.910 77.750 35.240 77.780 ;
        RECT 34.540 77.565 35.240 77.750 ;
        RECT 34.910 77.540 35.240 77.565 ;
        RECT 27.760 76.775 28.090 77.405 ;
        RECT 27.040 76.435 28.420 76.605 ;
        RECT 34.910 76.550 35.140 77.370 ;
        RECT 35.410 77.350 35.640 77.830 ;
        RECT 41.905 77.750 42.235 77.780 ;
        RECT 41.535 77.565 42.235 77.750 ;
        RECT 41.905 77.540 42.235 77.565 ;
        RECT 35.310 76.720 35.640 77.350 ;
        RECT 41.905 76.550 42.135 77.370 ;
        RECT 42.405 77.350 42.635 77.830 ;
        RECT 42.305 76.720 42.635 77.350 ;
        RECT 34.590 76.380 35.970 76.550 ;
        RECT 41.585 76.380 42.965 76.550 ;
        RECT 21.690 76.280 22.365 76.340 ;
        RECT 20.110 76.170 22.365 76.280 ;
        RECT 20.110 76.110 21.860 76.170 ;
        RECT 58.750 70.540 60.700 70.710 ;
        RECT 58.750 68.205 58.920 70.540 ;
        RECT 59.550 70.030 59.900 70.200 ;
        RECT 57.100 68.035 58.925 68.205 ;
        RECT 57.440 66.895 57.650 68.035 ;
        RECT 58.320 68.030 58.925 68.035 ;
        RECT 57.820 66.945 58.150 67.865 ;
        RECT 58.750 67.050 58.920 68.030 ;
        RECT 59.320 67.775 59.490 69.815 ;
        RECT 59.960 67.775 60.130 69.815 ;
        RECT 59.550 67.390 59.900 67.560 ;
        RECT 60.530 67.050 60.700 70.540 ;
        RECT 57.820 66.885 58.565 66.945 ;
        RECT 57.920 66.775 58.565 66.885 ;
        RECT 58.750 66.880 60.700 67.050 ;
        RECT 57.420 66.660 57.750 66.715 ;
        RECT 56.960 66.480 57.750 66.660 ;
        RECT 57.420 66.475 57.750 66.480 ;
        RECT 57.420 65.485 57.650 66.305 ;
        RECT 57.920 66.285 58.150 66.775 ;
        RECT 57.820 65.655 58.150 66.285 ;
        RECT 58.860 66.280 60.610 66.450 ;
        RECT 58.860 65.500 59.030 66.280 ;
        RECT 59.570 65.770 59.900 65.940 ;
        RECT 58.320 65.485 59.035 65.500 ;
        RECT 57.100 65.325 59.035 65.485 ;
        RECT 57.100 65.315 58.480 65.325 ;
        RECT 58.860 64.460 59.030 65.325 ;
        RECT 59.430 65.140 59.600 65.600 ;
        RECT 59.870 65.140 60.040 65.600 ;
        RECT 59.570 64.800 59.900 64.970 ;
        RECT 60.440 64.460 60.610 66.280 ;
        RECT 58.860 64.290 60.610 64.460 ;
        RECT 58.620 41.045 60.570 41.215 ;
        RECT 58.620 38.710 58.790 41.045 ;
        RECT 59.420 40.535 59.770 40.705 ;
        RECT 56.970 38.540 58.795 38.710 ;
        RECT 57.310 37.400 57.520 38.540 ;
        RECT 58.190 38.535 58.795 38.540 ;
        RECT 57.690 37.450 58.020 38.370 ;
        RECT 58.620 37.555 58.790 38.535 ;
        RECT 59.190 38.280 59.360 40.320 ;
        RECT 59.830 38.280 60.000 40.320 ;
        RECT 59.420 37.895 59.770 38.065 ;
        RECT 60.400 37.555 60.570 41.045 ;
        RECT 57.690 37.390 58.435 37.450 ;
        RECT 57.790 37.280 58.435 37.390 ;
        RECT 58.620 37.385 60.570 37.555 ;
        RECT 57.290 37.165 57.620 37.220 ;
        RECT 56.830 36.985 57.620 37.165 ;
        RECT 57.290 36.980 57.620 36.985 ;
        RECT 57.290 35.990 57.520 36.810 ;
        RECT 57.790 36.790 58.020 37.280 ;
        RECT 57.690 36.160 58.020 36.790 ;
        RECT 58.730 36.785 60.480 36.955 ;
        RECT 58.730 36.005 58.900 36.785 ;
        RECT 59.440 36.275 59.770 36.445 ;
        RECT 58.190 35.990 58.905 36.005 ;
        RECT 56.970 35.830 58.905 35.990 ;
        RECT 56.970 35.820 58.350 35.830 ;
        RECT 58.730 34.965 58.900 35.830 ;
        RECT 59.300 35.645 59.470 36.105 ;
        RECT 59.740 35.645 59.910 36.105 ;
        RECT 59.440 35.305 59.770 35.475 ;
        RECT 60.310 34.965 60.480 36.785 ;
        RECT 58.730 34.795 60.480 34.965 ;
        RECT 59.650 9.330 61.600 9.500 ;
        RECT 59.650 6.995 59.820 9.330 ;
        RECT 60.450 8.820 60.800 8.990 ;
        RECT 58.000 6.825 59.825 6.995 ;
        RECT 58.340 5.685 58.550 6.825 ;
        RECT 59.220 6.820 59.825 6.825 ;
        RECT 58.720 5.735 59.050 6.655 ;
        RECT 59.650 5.840 59.820 6.820 ;
        RECT 60.220 6.565 60.390 8.605 ;
        RECT 60.860 6.565 61.030 8.605 ;
        RECT 60.450 6.180 60.800 6.350 ;
        RECT 61.430 5.840 61.600 9.330 ;
        RECT 58.720 5.675 59.465 5.735 ;
        RECT 58.820 5.565 59.465 5.675 ;
        RECT 59.650 5.670 61.600 5.840 ;
        RECT 58.320 5.450 58.650 5.505 ;
        RECT 57.860 5.270 58.650 5.450 ;
        RECT 58.320 5.265 58.650 5.270 ;
        RECT 58.320 4.275 58.550 5.095 ;
        RECT 58.820 5.075 59.050 5.565 ;
        RECT 58.720 4.445 59.050 5.075 ;
        RECT 59.760 5.070 61.510 5.240 ;
        RECT 59.760 4.290 59.930 5.070 ;
        RECT 60.470 4.560 60.800 4.730 ;
        RECT 59.220 4.275 59.935 4.290 ;
        RECT 58.000 4.115 59.935 4.275 ;
        RECT 58.000 4.105 59.380 4.115 ;
        RECT 59.760 3.250 59.930 4.115 ;
        RECT 60.330 3.930 60.500 4.390 ;
        RECT 60.770 3.930 60.940 4.390 ;
        RECT 60.470 3.590 60.800 3.760 ;
        RECT 61.340 3.250 61.510 5.070 ;
        RECT 59.760 3.080 61.510 3.250 ;
      LAYER met1 ;
        RECT 58.350 222.450 58.650 222.480 ;
        RECT 56.050 222.150 58.650 222.450 ;
        RECT 47.950 219.450 48.250 219.480 ;
        RECT 51.350 219.450 51.650 219.480 ;
        RECT 47.950 219.150 51.650 219.450 ;
        RECT 47.950 219.120 48.250 219.150 ;
        RECT 51.350 219.120 51.650 219.150 ;
        RECT 56.050 213.920 56.350 222.150 ;
        RECT 58.350 222.120 58.650 222.150 ;
        RECT 55.250 213.150 55.550 213.180 ;
        RECT 47.120 212.850 55.550 213.150 ;
        RECT 55.250 212.820 55.550 212.850 ;
        RECT 54.250 212.050 54.550 212.080 ;
        RECT 47.120 211.750 54.550 212.050 ;
        RECT 54.250 211.720 54.550 211.750 ;
        RECT 16.620 208.440 16.940 208.500 ;
        RECT 17.540 208.440 17.860 208.500 ;
        RECT 16.620 208.300 17.860 208.440 ;
        RECT 16.620 208.240 16.940 208.300 ;
        RECT 17.540 208.240 17.860 208.300 ;
        RECT 25.820 208.100 26.140 208.160 ;
        RECT 29.040 208.100 29.360 208.160 ;
        RECT 25.820 207.960 29.360 208.100 ;
        RECT 25.820 207.900 26.140 207.960 ;
        RECT 29.040 207.900 29.360 207.960 ;
        RECT 8.270 207.280 43.230 207.760 ;
        RECT 17.540 206.880 17.860 207.140 ;
        RECT 22.600 207.080 22.920 207.140 ;
        RECT 30.420 207.080 30.740 207.140 ;
        RECT 20.850 206.940 30.740 207.080 ;
        RECT 14.795 206.740 15.085 206.785 ;
        RECT 17.080 206.740 17.400 206.800 ;
        RECT 14.795 206.600 17.400 206.740 ;
        RECT 14.795 206.555 15.085 206.600 ;
        RECT 17.080 206.540 17.400 206.600 ;
        RECT 11.100 206.400 11.420 206.460 ;
        RECT 11.575 206.400 11.865 206.445 ;
        RECT 11.100 206.260 11.865 206.400 ;
        RECT 11.100 206.200 11.420 206.260 ;
        RECT 11.575 206.215 11.865 206.260 ;
        RECT 12.955 206.400 13.245 206.445 ;
        RECT 13.860 206.400 14.180 206.460 ;
        RECT 12.955 206.260 14.180 206.400 ;
        RECT 12.955 206.215 13.245 206.260 ;
        RECT 13.860 206.200 14.180 206.260 ;
        RECT 18.000 206.200 18.320 206.460 ;
        RECT 20.850 206.445 20.990 206.940 ;
        RECT 22.600 206.880 22.920 206.940 ;
        RECT 30.420 206.880 30.740 206.940 ;
        RECT 31.800 207.080 32.120 207.140 ;
        RECT 35.495 207.080 35.785 207.125 ;
        RECT 31.800 206.940 35.785 207.080 ;
        RECT 31.800 206.880 32.120 206.940 ;
        RECT 35.495 206.895 35.785 206.940 ;
        RECT 38.240 206.880 38.560 207.140 ;
        RECT 40.555 207.080 40.845 207.125 ;
        RECT 47.900 207.080 48.220 207.140 ;
        RECT 40.555 206.940 48.220 207.080 ;
        RECT 40.555 206.895 40.845 206.940 ;
        RECT 47.900 206.880 48.220 206.940 ;
        RECT 26.295 206.740 26.585 206.785 ;
        RECT 23.610 206.600 26.585 206.740 ;
        RECT 23.610 206.460 23.750 206.600 ;
        RECT 26.295 206.555 26.585 206.600 ;
        RECT 26.755 206.740 27.045 206.785 ;
        RECT 29.040 206.740 29.360 206.800 ;
        RECT 34.560 206.740 34.880 206.800 ;
        RECT 26.755 206.600 28.350 206.740 ;
        RECT 26.755 206.555 27.045 206.600 ;
        RECT 28.210 206.460 28.350 206.600 ;
        RECT 29.040 206.600 34.880 206.740 ;
        RECT 29.040 206.540 29.360 206.600 ;
        RECT 34.560 206.540 34.880 206.600 ;
        RECT 19.855 206.400 20.145 206.445 ;
        RECT 18.550 206.260 20.145 206.400 ;
        RECT 18.550 205.780 18.690 206.260 ;
        RECT 19.855 206.215 20.145 206.260 ;
        RECT 20.775 206.215 21.065 206.445 ;
        RECT 23.520 206.200 23.840 206.460 ;
        RECT 24.455 206.215 24.745 206.445 ;
        RECT 25.375 206.400 25.665 206.445 ;
        RECT 25.820 206.400 26.140 206.460 ;
        RECT 25.375 206.260 26.140 206.400 ;
        RECT 25.375 206.215 25.665 206.260 ;
        RECT 22.140 206.060 22.460 206.120 ;
        RECT 23.075 206.060 23.365 206.105 ;
        RECT 22.140 205.920 23.365 206.060 ;
        RECT 24.530 206.060 24.670 206.215 ;
        RECT 25.820 206.200 26.140 206.260 ;
        RECT 27.215 206.400 27.505 206.445 ;
        RECT 27.660 206.400 27.980 206.460 ;
        RECT 27.215 206.260 27.980 206.400 ;
        RECT 27.215 206.215 27.505 206.260 ;
        RECT 27.660 206.200 27.980 206.260 ;
        RECT 28.120 206.200 28.440 206.460 ;
        RECT 29.130 206.400 29.270 206.540 ;
        RECT 29.515 206.400 29.805 206.445 ;
        RECT 31.340 206.400 31.660 206.460 ;
        RECT 35.035 206.400 35.325 206.445 ;
        RECT 29.130 206.260 29.805 206.400 ;
        RECT 29.515 206.215 29.805 206.260 ;
        RECT 30.050 206.260 31.110 206.400 ;
        RECT 30.050 206.060 30.190 206.260 ;
        RECT 24.530 205.920 30.190 206.060 ;
        RECT 22.140 205.860 22.460 205.920 ;
        RECT 23.075 205.875 23.365 205.920 ;
        RECT 30.420 205.860 30.740 206.120 ;
        RECT 30.970 206.060 31.110 206.260 ;
        RECT 31.340 206.260 35.325 206.400 ;
        RECT 31.340 206.200 31.660 206.260 ;
        RECT 35.035 206.215 35.325 206.260 ;
        RECT 36.860 206.400 37.180 206.460 ;
        RECT 37.335 206.400 37.625 206.445 ;
        RECT 36.860 206.260 37.625 206.400 ;
        RECT 36.860 206.200 37.180 206.260 ;
        RECT 37.335 206.215 37.625 206.260 ;
        RECT 40.540 206.400 40.860 206.460 ;
        RECT 41.015 206.400 41.305 206.445 ;
        RECT 40.540 206.260 41.305 206.400 ;
        RECT 40.540 206.200 40.860 206.260 ;
        RECT 41.015 206.215 41.305 206.260 ;
        RECT 35.480 206.060 35.800 206.120 ;
        RECT 30.970 205.920 35.800 206.060 ;
        RECT 35.480 205.860 35.800 205.920 ;
        RECT 10.195 205.535 10.485 205.765 ;
        RECT 6.040 205.380 6.360 205.440 ;
        RECT 10.270 205.380 10.410 205.535 ;
        RECT 18.460 205.520 18.780 205.780 ;
        RECT 28.135 205.720 28.425 205.765 ;
        RECT 34.100 205.720 34.420 205.780 ;
        RECT 28.135 205.580 34.420 205.720 ;
        RECT 28.135 205.535 28.425 205.580 ;
        RECT 34.100 205.520 34.420 205.580 ;
        RECT 6.040 205.240 10.410 205.380 ;
        RECT 15.240 205.380 15.560 205.440 ;
        RECT 18.935 205.380 19.225 205.425 ;
        RECT 15.240 205.240 19.225 205.380 ;
        RECT 6.040 205.180 6.360 205.240 ;
        RECT 15.240 205.180 15.560 205.240 ;
        RECT 18.935 205.195 19.225 205.240 ;
        RECT 28.580 205.180 28.900 205.440 ;
        RECT 8.270 204.560 43.230 205.040 ;
        RECT 10.180 204.160 10.500 204.420 ;
        RECT 12.495 204.360 12.785 204.405 ;
        RECT 13.860 204.360 14.180 204.420 ;
        RECT 12.495 204.220 14.180 204.360 ;
        RECT 12.495 204.175 12.785 204.220 ;
        RECT 13.860 204.160 14.180 204.220 ;
        RECT 14.780 204.360 15.100 204.420 ;
        RECT 27.675 204.360 27.965 204.405 ;
        RECT 14.780 204.220 27.965 204.360 ;
        RECT 14.780 204.160 15.100 204.220 ;
        RECT 27.675 204.175 27.965 204.220 ;
        RECT 34.100 204.360 34.420 204.420 ;
        RECT 34.100 204.220 36.630 204.360 ;
        RECT 18.015 204.020 18.305 204.065 ;
        RECT 26.740 204.020 27.060 204.080 ;
        RECT 10.270 203.880 16.390 204.020 ;
        RECT 10.270 203.060 10.410 203.880 ;
        RECT 15.240 203.680 15.560 203.740 ;
        RECT 13.490 203.540 15.560 203.680 ;
        RECT 11.100 203.140 11.420 203.400 ;
        RECT 13.490 203.385 13.630 203.540 ;
        RECT 15.240 203.480 15.560 203.540 ;
        RECT 16.250 203.400 16.390 203.880 ;
        RECT 18.015 203.880 27.060 204.020 ;
        RECT 18.015 203.835 18.305 203.880 ;
        RECT 26.740 203.820 27.060 203.880 ;
        RECT 27.750 203.680 27.890 204.175 ;
        RECT 34.100 204.160 34.420 204.220 ;
        RECT 30.535 204.020 30.825 204.065 ;
        RECT 33.655 204.020 33.945 204.065 ;
        RECT 35.545 204.020 35.835 204.065 ;
        RECT 30.535 203.880 35.835 204.020 ;
        RECT 36.490 204.020 36.630 204.220 ;
        RECT 36.860 204.160 37.180 204.420 ;
        RECT 36.490 203.880 40.310 204.020 ;
        RECT 30.535 203.835 30.825 203.880 ;
        RECT 33.655 203.835 33.945 203.880 ;
        RECT 35.545 203.835 35.835 203.880 ;
        RECT 37.320 203.680 37.640 203.740 ;
        RECT 23.150 203.540 26.050 203.680 ;
        RECT 27.750 203.540 38.010 203.680 ;
        RECT 13.415 203.155 13.705 203.385 ;
        RECT 13.860 203.340 14.180 203.400 ;
        RECT 14.780 203.340 15.100 203.400 ;
        RECT 13.860 203.200 15.100 203.340 ;
        RECT 13.860 203.140 14.180 203.200 ;
        RECT 14.780 203.140 15.100 203.200 ;
        RECT 15.715 203.320 16.005 203.385 ;
        RECT 16.160 203.320 16.480 203.400 ;
        RECT 15.715 203.180 16.480 203.320 ;
        RECT 15.715 203.155 16.005 203.180 ;
        RECT 16.160 203.140 16.480 203.180 ;
        RECT 16.635 203.340 16.925 203.385 ;
        RECT 23.150 203.340 23.290 203.540 ;
        RECT 25.910 203.400 26.050 203.540 ;
        RECT 37.320 203.480 37.640 203.540 ;
        RECT 16.635 203.200 23.290 203.340 ;
        RECT 23.520 203.340 23.840 203.400 ;
        RECT 24.455 203.340 24.745 203.385 ;
        RECT 23.520 203.200 24.745 203.340 ;
        RECT 16.635 203.155 16.925 203.200 ;
        RECT 10.180 202.800 10.500 203.060 ;
        RECT 11.190 202.660 11.330 203.140 ;
        RECT 11.560 202.800 11.880 203.060 ;
        RECT 15.255 203.000 15.545 203.045 ;
        RECT 17.080 203.000 17.400 203.060 ;
        RECT 15.255 202.860 17.400 203.000 ;
        RECT 15.255 202.815 15.545 202.860 ;
        RECT 17.080 202.800 17.400 202.860 ;
        RECT 13.875 202.660 14.165 202.705 ;
        RECT 11.190 202.520 14.165 202.660 ;
        RECT 13.875 202.475 14.165 202.520 ;
        RECT 14.320 202.660 14.640 202.720 ;
        RECT 17.630 202.660 17.770 203.200 ;
        RECT 23.520 203.140 23.840 203.200 ;
        RECT 24.455 203.155 24.745 203.200 ;
        RECT 25.820 203.140 26.140 203.400 ;
        RECT 26.280 203.340 26.600 203.400 ;
        RECT 29.455 203.340 29.745 203.360 ;
        RECT 26.280 203.200 29.745 203.340 ;
        RECT 26.280 203.140 26.600 203.200 ;
        RECT 29.455 203.045 29.745 203.200 ;
        RECT 30.535 203.340 30.825 203.385 ;
        RECT 34.115 203.340 34.405 203.385 ;
        RECT 35.950 203.340 36.240 203.385 ;
        RECT 30.535 203.200 36.240 203.340 ;
        RECT 30.535 203.155 30.825 203.200 ;
        RECT 34.115 203.155 34.405 203.200 ;
        RECT 35.950 203.155 36.240 203.200 ;
        RECT 36.400 203.140 36.720 203.400 ;
        RECT 37.870 203.385 38.010 203.540 ;
        RECT 40.170 203.385 40.310 203.880 ;
        RECT 37.795 203.155 38.085 203.385 ;
        RECT 39.635 203.155 39.925 203.385 ;
        RECT 40.095 203.155 40.385 203.385 ;
        RECT 18.935 203.000 19.225 203.045 ;
        RECT 29.155 203.000 29.745 203.045 ;
        RECT 32.395 203.000 33.045 203.045 ;
        RECT 18.935 202.860 28.810 203.000 ;
        RECT 18.935 202.815 19.225 202.860 ;
        RECT 14.320 202.520 17.770 202.660 ;
        RECT 19.380 202.660 19.700 202.720 ;
        RECT 21.695 202.660 21.985 202.705 ;
        RECT 19.380 202.520 21.985 202.660 ;
        RECT 28.670 202.660 28.810 202.860 ;
        RECT 29.155 202.860 33.045 203.000 ;
        RECT 29.155 202.815 29.445 202.860 ;
        RECT 32.395 202.815 33.045 202.860 ;
        RECT 35.020 202.800 35.340 203.060 ;
        RECT 38.240 202.800 38.560 203.060 ;
        RECT 38.715 202.815 39.005 203.045 ;
        RECT 39.710 203.000 39.850 203.155 ;
        RECT 43.760 203.140 44.080 203.400 ;
        RECT 43.850 203.000 43.990 203.140 ;
        RECT 39.710 202.860 43.990 203.000 ;
        RECT 30.420 202.660 30.740 202.720 ;
        RECT 28.670 202.520 30.740 202.660 ;
        RECT 14.320 202.460 14.640 202.520 ;
        RECT 19.380 202.460 19.700 202.520 ;
        RECT 21.695 202.475 21.985 202.520 ;
        RECT 30.420 202.460 30.740 202.520 ;
        RECT 31.800 202.660 32.120 202.720 ;
        RECT 38.790 202.660 38.930 202.815 ;
        RECT 31.800 202.520 38.930 202.660 ;
        RECT 41.015 202.660 41.305 202.705 ;
        RECT 43.300 202.660 43.620 202.720 ;
        RECT 41.015 202.520 43.620 202.660 ;
        RECT 31.800 202.460 32.120 202.520 ;
        RECT 41.015 202.475 41.305 202.520 ;
        RECT 43.300 202.460 43.620 202.520 ;
        RECT 8.270 201.840 43.230 202.320 ;
        RECT 11.115 201.640 11.405 201.685 ;
        RECT 11.560 201.640 11.880 201.700 ;
        RECT 11.115 201.500 11.880 201.640 ;
        RECT 11.115 201.455 11.405 201.500 ;
        RECT 11.560 201.440 11.880 201.500 ;
        RECT 14.335 201.640 14.625 201.685 ;
        RECT 14.780 201.640 15.100 201.700 ;
        RECT 23.520 201.640 23.840 201.700 ;
        RECT 14.335 201.500 23.840 201.640 ;
        RECT 14.335 201.455 14.625 201.500 ;
        RECT 14.780 201.440 15.100 201.500 ;
        RECT 23.520 201.440 23.840 201.500 ;
        RECT 28.580 201.440 28.900 201.700 ;
        RECT 33.195 201.640 33.485 201.685 ;
        RECT 35.020 201.640 35.340 201.700 ;
        RECT 33.195 201.500 35.340 201.640 ;
        RECT 33.195 201.455 33.485 201.500 ;
        RECT 35.020 201.440 35.340 201.500 ;
        RECT 35.480 201.640 35.800 201.700 ;
        RECT 38.255 201.640 38.545 201.685 ;
        RECT 35.480 201.500 38.545 201.640 ;
        RECT 35.480 201.440 35.800 201.500 ;
        RECT 38.255 201.455 38.545 201.500 ;
        RECT 12.955 201.300 13.245 201.345 ;
        RECT 15.815 201.300 16.105 201.345 ;
        RECT 19.055 201.300 19.705 201.345 ;
        RECT 21.220 201.300 21.540 201.360 ;
        RECT 26.280 201.300 26.600 201.360 ;
        RECT 11.190 201.160 15.470 201.300 ;
        RECT 11.190 201.020 11.330 201.160 ;
        RECT 12.955 201.115 13.245 201.160 ;
        RECT 9.720 200.760 10.040 201.020 ;
        RECT 11.100 200.760 11.420 201.020 ;
        RECT 12.035 200.775 12.325 201.005 ;
        RECT 13.415 200.960 13.705 201.005 ;
        RECT 14.320 200.960 14.640 201.020 ;
        RECT 13.415 200.820 14.640 200.960 ;
        RECT 15.330 200.960 15.470 201.160 ;
        RECT 15.815 201.160 26.600 201.300 ;
        RECT 15.815 201.115 16.405 201.160 ;
        RECT 19.055 201.115 19.705 201.160 ;
        RECT 15.330 200.820 15.930 200.960 ;
        RECT 13.415 200.775 13.705 200.820 ;
        RECT 12.110 200.620 12.250 200.775 ;
        RECT 14.320 200.760 14.640 200.820 ;
        RECT 15.240 200.620 15.560 200.680 ;
        RECT 12.110 200.480 15.560 200.620 ;
        RECT 15.790 200.620 15.930 200.820 ;
        RECT 16.115 200.800 16.405 201.115 ;
        RECT 21.220 201.100 21.540 201.160 ;
        RECT 26.280 201.100 26.600 201.160 ;
        RECT 17.195 200.960 17.485 201.005 ;
        RECT 20.775 200.960 21.065 201.005 ;
        RECT 22.610 200.960 22.900 201.005 ;
        RECT 17.195 200.820 22.900 200.960 ;
        RECT 17.195 200.775 17.485 200.820 ;
        RECT 20.775 200.775 21.065 200.820 ;
        RECT 22.610 200.775 22.900 200.820 ;
        RECT 23.060 200.760 23.380 201.020 ;
        RECT 24.915 200.960 25.205 201.005 ;
        RECT 28.670 200.960 28.810 201.440 ;
        RECT 30.420 201.300 30.740 201.360 ;
        RECT 30.420 201.160 35.710 201.300 ;
        RECT 30.420 201.100 30.740 201.160 ;
        RECT 35.570 201.020 35.710 201.160 ;
        RECT 36.030 201.160 41.230 201.300 ;
        RECT 36.030 201.020 36.170 201.160 ;
        RECT 24.915 200.820 28.810 200.960 ;
        RECT 29.040 200.960 29.360 201.020 ;
        RECT 31.800 200.960 32.120 201.020 ;
        RECT 29.040 200.820 32.120 200.960 ;
        RECT 24.915 200.775 25.205 200.820 ;
        RECT 29.040 200.760 29.360 200.820 ;
        RECT 31.800 200.760 32.120 200.820 ;
        RECT 34.560 200.760 34.880 201.020 ;
        RECT 35.480 200.760 35.800 201.020 ;
        RECT 35.940 200.760 36.260 201.020 ;
        RECT 37.320 200.760 37.640 201.020 ;
        RECT 37.780 200.960 38.100 201.020 ;
        RECT 39.175 200.960 39.465 201.005 ;
        RECT 37.780 200.820 39.465 200.960 ;
        RECT 37.780 200.760 38.100 200.820 ;
        RECT 39.175 200.775 39.465 200.820 ;
        RECT 39.635 200.775 39.925 201.005 ;
        RECT 18.920 200.620 19.240 200.680 ;
        RECT 21.220 200.620 21.540 200.680 ;
        RECT 15.790 200.480 16.620 200.620 ;
        RECT 15.240 200.420 15.560 200.480 ;
        RECT 10.640 199.740 10.960 200.000 ;
        RECT 16.480 199.940 16.620 200.480 ;
        RECT 18.920 200.480 21.540 200.620 ;
        RECT 18.920 200.420 19.240 200.480 ;
        RECT 21.220 200.420 21.540 200.480 ;
        RECT 21.695 200.620 21.985 200.665 ;
        RECT 26.295 200.620 26.585 200.665 ;
        RECT 21.695 200.480 26.585 200.620 ;
        RECT 21.695 200.435 21.985 200.480 ;
        RECT 26.295 200.435 26.585 200.480 ;
        RECT 27.660 200.620 27.980 200.680 ;
        RECT 28.580 200.620 28.900 200.680 ;
        RECT 29.975 200.620 30.265 200.665 ;
        RECT 27.660 200.480 30.265 200.620 ;
        RECT 34.650 200.620 34.790 200.760 ;
        RECT 39.710 200.620 39.850 200.775 ;
        RECT 40.080 200.760 40.400 201.020 ;
        RECT 41.090 201.005 41.230 201.160 ;
        RECT 41.015 200.775 41.305 201.005 ;
        RECT 34.650 200.480 39.850 200.620 ;
        RECT 27.660 200.420 27.980 200.480 ;
        RECT 28.580 200.420 28.900 200.480 ;
        RECT 29.975 200.435 30.265 200.480 ;
        RECT 17.195 200.280 17.485 200.325 ;
        RECT 20.315 200.280 20.605 200.325 ;
        RECT 22.205 200.280 22.495 200.325 ;
        RECT 17.195 200.140 22.495 200.280 ;
        RECT 17.195 200.095 17.485 200.140 ;
        RECT 20.315 200.095 20.605 200.140 ;
        RECT 22.205 200.095 22.495 200.140 ;
        RECT 25.835 200.280 26.125 200.325 ;
        RECT 31.340 200.280 31.660 200.340 ;
        RECT 25.835 200.140 31.660 200.280 ;
        RECT 25.835 200.095 26.125 200.140 ;
        RECT 31.340 200.080 31.660 200.140 ;
        RECT 22.600 199.940 22.920 200.000 ;
        RECT 16.480 199.800 22.920 199.940 ;
        RECT 22.600 199.740 22.920 199.800 ;
        RECT 32.260 199.940 32.580 200.000 ;
        RECT 34.575 199.940 34.865 199.985 ;
        RECT 32.260 199.800 34.865 199.940 ;
        RECT 32.260 199.740 32.580 199.800 ;
        RECT 34.575 199.755 34.865 199.800 ;
        RECT 35.020 199.940 35.340 200.000 ;
        RECT 38.240 199.940 38.560 200.000 ;
        RECT 35.020 199.800 38.560 199.940 ;
        RECT 35.020 199.740 35.340 199.800 ;
        RECT 38.240 199.740 38.560 199.800 ;
        RECT 8.270 199.120 43.230 199.600 ;
        RECT 11.560 198.920 11.880 198.980 ;
        RECT 14.320 198.920 14.640 198.980 ;
        RECT 10.270 198.780 11.330 198.920 ;
        RECT 7.420 198.240 7.740 198.300 ;
        RECT 10.270 198.240 10.410 198.780 ;
        RECT 10.640 198.380 10.960 198.640 ;
        RECT 11.190 198.625 11.330 198.780 ;
        RECT 11.560 198.780 14.640 198.920 ;
        RECT 11.560 198.720 11.880 198.780 ;
        RECT 14.320 198.720 14.640 198.780 ;
        RECT 30.895 198.920 31.185 198.965 ;
        RECT 31.800 198.920 32.120 198.980 ;
        RECT 30.895 198.780 40.310 198.920 ;
        RECT 30.895 198.735 31.185 198.780 ;
        RECT 31.800 198.720 32.120 198.780 ;
        RECT 11.115 198.395 11.405 198.625 ;
        RECT 18.460 198.580 18.780 198.640 ;
        RECT 33.755 198.580 34.045 198.625 ;
        RECT 36.875 198.580 37.165 198.625 ;
        RECT 38.765 198.580 39.055 198.625 ;
        RECT 15.790 198.440 23.980 198.580 ;
        RECT 7.420 198.100 10.410 198.240 ;
        RECT 7.420 198.040 7.740 198.100 ;
        RECT 10.195 197.900 10.485 197.945 ;
        RECT 10.730 197.900 10.870 198.380 ;
        RECT 10.195 197.760 10.870 197.900 ;
        RECT 10.195 197.715 10.485 197.760 ;
        RECT 14.780 197.700 15.100 197.960 ;
        RECT 15.240 197.945 15.560 197.960 ;
        RECT 15.240 197.900 15.645 197.945 ;
        RECT 15.790 197.900 15.930 198.440 ;
        RECT 18.460 198.380 18.780 198.440 ;
        RECT 16.160 198.040 16.480 198.300 ;
        RECT 18.935 198.240 19.225 198.285 ;
        RECT 19.840 198.240 20.160 198.300 ;
        RECT 18.935 198.100 20.160 198.240 ;
        RECT 18.935 198.055 19.225 198.100 ;
        RECT 19.840 198.040 20.160 198.100 ;
        RECT 20.300 198.240 20.620 198.300 ;
        RECT 23.840 198.240 23.980 198.440 ;
        RECT 33.755 198.440 39.055 198.580 ;
        RECT 33.755 198.395 34.045 198.440 ;
        RECT 36.875 198.395 37.165 198.440 ;
        RECT 38.765 198.395 39.055 198.440 ;
        RECT 40.170 198.300 40.310 198.780 ;
        RECT 29.500 198.240 29.820 198.300 ;
        RECT 35.940 198.240 36.260 198.300 ;
        RECT 20.300 198.100 22.830 198.240 ;
        RECT 23.840 198.100 29.820 198.240 ;
        RECT 20.300 198.040 20.620 198.100 ;
        RECT 15.240 197.760 15.930 197.900 ;
        RECT 16.250 197.900 16.390 198.040 ;
        RECT 16.635 197.900 16.925 197.945 ;
        RECT 16.250 197.760 16.925 197.900 ;
        RECT 15.240 197.715 15.645 197.760 ;
        RECT 16.635 197.715 16.925 197.760 ;
        RECT 17.095 197.900 17.385 197.945 ;
        RECT 17.540 197.900 17.860 197.960 ;
        RECT 22.690 197.945 22.830 198.100 ;
        RECT 24.070 197.945 24.210 198.100 ;
        RECT 29.500 198.040 29.820 198.100 ;
        RECT 31.890 198.100 36.260 198.240 ;
        RECT 17.095 197.760 17.860 197.900 ;
        RECT 17.095 197.715 17.385 197.760 ;
        RECT 15.240 197.700 15.560 197.715 ;
        RECT 17.540 197.700 17.860 197.760 ;
        RECT 22.615 197.715 22.905 197.945 ;
        RECT 23.995 197.715 24.285 197.945 ;
        RECT 27.200 197.900 27.520 197.960 ;
        RECT 29.975 197.900 30.265 197.945 ;
        RECT 27.200 197.760 30.265 197.900 ;
        RECT 14.335 197.560 14.625 197.605 ;
        RECT 10.730 197.420 14.625 197.560 ;
        RECT 14.870 197.560 15.010 197.700 ;
        RECT 16.175 197.560 16.465 197.605 ;
        RECT 14.870 197.420 16.465 197.560 ;
        RECT 10.180 197.220 10.500 197.280 ;
        RECT 10.730 197.220 10.870 197.420 ;
        RECT 14.335 197.375 14.625 197.420 ;
        RECT 16.175 197.375 16.465 197.420 ;
        RECT 20.315 197.560 20.605 197.605 ;
        RECT 21.695 197.560 21.985 197.605 ;
        RECT 20.315 197.420 21.985 197.560 ;
        RECT 22.690 197.560 22.830 197.715 ;
        RECT 27.200 197.700 27.520 197.760 ;
        RECT 29.975 197.715 30.265 197.760 ;
        RECT 28.120 197.560 28.440 197.620 ;
        RECT 31.890 197.560 32.030 198.100 ;
        RECT 35.940 198.040 36.260 198.100 ;
        RECT 36.400 198.240 36.720 198.300 ;
        RECT 39.635 198.240 39.925 198.285 ;
        RECT 36.400 198.100 39.925 198.240 ;
        RECT 36.400 198.040 36.720 198.100 ;
        RECT 39.635 198.055 39.925 198.100 ;
        RECT 40.080 198.040 40.400 198.300 ;
        RECT 32.675 197.605 32.965 197.920 ;
        RECT 33.755 197.900 34.045 197.945 ;
        RECT 37.335 197.900 37.625 197.945 ;
        RECT 39.170 197.900 39.460 197.945 ;
        RECT 33.755 197.760 39.460 197.900 ;
        RECT 33.755 197.715 34.045 197.760 ;
        RECT 37.335 197.715 37.625 197.760 ;
        RECT 39.170 197.715 39.460 197.760 ;
        RECT 22.690 197.420 32.030 197.560 ;
        RECT 32.375 197.560 32.965 197.605 ;
        RECT 35.615 197.560 36.265 197.605 ;
        RECT 32.375 197.420 36.265 197.560 ;
        RECT 20.315 197.375 20.605 197.420 ;
        RECT 21.695 197.375 21.985 197.420 ;
        RECT 28.120 197.360 28.440 197.420 ;
        RECT 32.375 197.375 32.665 197.420 ;
        RECT 10.180 197.080 10.870 197.220 ;
        RECT 10.180 197.020 10.500 197.080 ;
        RECT 13.860 197.020 14.180 197.280 ;
        RECT 18.000 197.020 18.320 197.280 ;
        RECT 22.600 197.220 22.920 197.280 ;
        RECT 23.535 197.220 23.825 197.265 ;
        RECT 27.660 197.220 27.980 197.280 ;
        RECT 22.600 197.080 27.980 197.220 ;
        RECT 22.600 197.020 22.920 197.080 ;
        RECT 23.535 197.035 23.825 197.080 ;
        RECT 27.660 197.020 27.980 197.080 ;
        RECT 29.055 197.220 29.345 197.265 ;
        RECT 30.880 197.220 31.200 197.280 ;
        RECT 29.055 197.080 31.200 197.220 ;
        RECT 29.055 197.035 29.345 197.080 ;
        RECT 30.880 197.020 31.200 197.080 ;
        RECT 31.800 197.220 32.120 197.280 ;
        RECT 32.810 197.220 32.950 197.420 ;
        RECT 35.615 197.375 36.265 197.420 ;
        RECT 38.255 197.560 38.545 197.605 ;
        RECT 38.700 197.560 39.020 197.620 ;
        RECT 38.255 197.420 39.020 197.560 ;
        RECT 38.255 197.375 38.545 197.420 ;
        RECT 38.700 197.360 39.020 197.420 ;
        RECT 31.800 197.080 32.950 197.220 ;
        RECT 31.800 197.020 32.120 197.080 ;
        RECT 8.270 196.400 43.230 196.880 ;
        RECT 9.720 196.000 10.040 196.260 ;
        RECT 17.080 196.200 17.400 196.260 ;
        RECT 20.300 196.200 20.620 196.260 ;
        RECT 10.730 196.060 20.620 196.200 ;
        RECT 10.730 195.565 10.870 196.060 ;
        RECT 17.080 196.000 17.400 196.060 ;
        RECT 20.300 196.000 20.620 196.060 ;
        RECT 21.005 196.200 21.295 196.245 ;
        RECT 22.600 196.200 22.920 196.260 ;
        RECT 21.005 196.060 22.920 196.200 ;
        RECT 21.005 196.015 21.295 196.060 ;
        RECT 22.600 196.000 22.920 196.060 ;
        RECT 35.110 196.060 40.310 196.200 ;
        RECT 18.920 195.905 19.240 195.920 ;
        RECT 12.960 195.860 13.250 195.905 ;
        RECT 14.820 195.860 15.110 195.905 ;
        RECT 12.960 195.720 15.110 195.860 ;
        RECT 12.960 195.675 13.250 195.720 ;
        RECT 14.820 195.675 15.110 195.720 ;
        RECT 15.740 195.860 16.030 195.905 ;
        RECT 18.920 195.860 19.290 195.905 ;
        RECT 23.060 195.860 23.380 195.920 ;
        RECT 15.740 195.720 19.290 195.860 ;
        RECT 15.740 195.675 16.030 195.720 ;
        RECT 18.920 195.675 19.290 195.720 ;
        RECT 21.770 195.720 23.380 195.860 ;
        RECT 10.655 195.520 10.945 195.565 ;
        RECT 9.350 195.380 10.945 195.520 ;
        RECT 9.350 194.900 9.490 195.380 ;
        RECT 10.655 195.335 10.945 195.380 ;
        RECT 11.100 195.320 11.420 195.580 ;
        RECT 14.895 195.520 15.110 195.675 ;
        RECT 18.920 195.660 19.240 195.675 ;
        RECT 17.140 195.520 17.430 195.565 ;
        RECT 12.110 195.380 14.550 195.520 ;
        RECT 14.895 195.380 17.430 195.520 ;
        RECT 12.110 195.225 12.250 195.380 ;
        RECT 12.035 194.995 12.325 195.225 ;
        RECT 13.860 194.980 14.180 195.240 ;
        RECT 14.410 195.180 14.550 195.380 ;
        RECT 17.140 195.335 17.430 195.380 ;
        RECT 16.620 195.180 16.940 195.240 ;
        RECT 21.770 195.225 21.910 195.720 ;
        RECT 23.060 195.660 23.380 195.720 ;
        RECT 25.355 195.860 26.005 195.905 ;
        RECT 26.280 195.860 26.600 195.920 ;
        RECT 28.955 195.860 29.245 195.905 ;
        RECT 25.355 195.720 29.245 195.860 ;
        RECT 25.355 195.675 26.005 195.720 ;
        RECT 26.280 195.660 26.600 195.720 ;
        RECT 28.655 195.675 29.245 195.720 ;
        RECT 29.590 195.720 34.790 195.860 ;
        RECT 22.160 195.520 22.450 195.565 ;
        RECT 23.995 195.520 24.285 195.565 ;
        RECT 27.575 195.520 27.865 195.565 ;
        RECT 22.160 195.380 27.865 195.520 ;
        RECT 22.160 195.335 22.450 195.380 ;
        RECT 23.995 195.335 24.285 195.380 ;
        RECT 27.575 195.335 27.865 195.380 ;
        RECT 28.655 195.360 28.945 195.675 ;
        RECT 29.590 195.580 29.730 195.720 ;
        RECT 34.650 195.580 34.790 195.720 ;
        RECT 35.110 195.580 35.250 196.060 ;
        RECT 35.495 195.860 35.785 195.905 ;
        RECT 38.240 195.860 38.560 195.920 ;
        RECT 35.495 195.720 38.560 195.860 ;
        RECT 35.495 195.675 35.785 195.720 ;
        RECT 38.240 195.660 38.560 195.720 ;
        RECT 39.620 195.660 39.940 195.920 ;
        RECT 29.500 195.320 29.820 195.580 ;
        RECT 31.815 195.335 32.105 195.565 ;
        RECT 21.695 195.180 21.985 195.225 ;
        RECT 14.410 195.040 21.985 195.180 ;
        RECT 16.620 194.980 16.940 195.040 ;
        RECT 21.695 194.995 21.985 195.040 ;
        RECT 23.060 194.980 23.380 195.240 ;
        RECT 25.820 195.180 26.140 195.240 ;
        RECT 31.890 195.180 32.030 195.335 ;
        RECT 34.560 195.320 34.880 195.580 ;
        RECT 35.020 195.520 35.340 195.580 ;
        RECT 35.955 195.520 36.245 195.565 ;
        RECT 35.020 195.380 36.245 195.520 ;
        RECT 35.020 195.320 35.340 195.380 ;
        RECT 35.955 195.335 36.245 195.380 ;
        RECT 36.415 195.335 36.705 195.565 ;
        RECT 36.860 195.520 37.180 195.580 ;
        RECT 38.715 195.520 39.005 195.565 ;
        RECT 36.860 195.380 39.005 195.520 ;
        RECT 25.820 195.040 32.030 195.180 ;
        RECT 25.820 194.980 26.140 195.040 ;
        RECT 9.260 194.640 9.580 194.900 ;
        RECT 12.500 194.840 12.790 194.885 ;
        RECT 14.360 194.840 14.650 194.885 ;
        RECT 17.140 194.840 17.430 194.885 ;
        RECT 12.500 194.700 17.430 194.840 ;
        RECT 12.500 194.655 12.790 194.700 ;
        RECT 14.360 194.655 14.650 194.700 ;
        RECT 17.140 194.655 17.430 194.700 ;
        RECT 18.000 194.840 18.320 194.900 ;
        RECT 22.565 194.840 22.855 194.885 ;
        RECT 24.455 194.840 24.745 194.885 ;
        RECT 27.575 194.840 27.865 194.885 ;
        RECT 18.000 194.700 22.370 194.840 ;
        RECT 18.000 194.640 18.320 194.700 ;
        RECT 13.860 194.500 14.180 194.560 ;
        RECT 19.380 194.500 19.700 194.560 ;
        RECT 13.860 194.360 19.700 194.500 ;
        RECT 22.230 194.500 22.370 194.700 ;
        RECT 22.565 194.700 27.865 194.840 ;
        RECT 22.565 194.655 22.855 194.700 ;
        RECT 24.455 194.655 24.745 194.700 ;
        RECT 27.575 194.655 27.865 194.700 ;
        RECT 35.940 194.840 36.260 194.900 ;
        RECT 36.490 194.840 36.630 195.335 ;
        RECT 36.860 195.320 37.180 195.380 ;
        RECT 38.715 195.335 39.005 195.380 ;
        RECT 39.175 195.335 39.465 195.565 ;
        RECT 40.170 195.520 40.310 196.060 ;
        RECT 40.555 195.520 40.845 195.565 ;
        RECT 40.170 195.380 40.845 195.520 ;
        RECT 40.555 195.335 40.845 195.380 ;
        RECT 38.240 195.180 38.560 195.240 ;
        RECT 39.250 195.180 39.390 195.335 ;
        RECT 43.760 195.180 44.080 195.240 ;
        RECT 38.240 195.040 44.080 195.180 ;
        RECT 53.250 195.050 53.550 195.080 ;
        RECT 38.240 194.980 38.560 195.040 ;
        RECT 43.760 194.980 44.080 195.040 ;
        RECT 36.860 194.840 37.180 194.900 ;
        RECT 35.940 194.700 37.180 194.840 ;
        RECT 35.940 194.640 36.260 194.700 ;
        RECT 36.860 194.640 37.180 194.700 ;
        RECT 37.335 194.840 37.625 194.885 ;
        RECT 41.920 194.840 42.240 194.900 ;
        RECT 37.335 194.700 42.240 194.840 ;
        RECT 47.520 194.750 53.550 195.050 ;
        RECT 53.250 194.720 53.550 194.750 ;
        RECT 37.335 194.655 37.625 194.700 ;
        RECT 41.920 194.640 42.240 194.700 ;
        RECT 28.580 194.500 28.900 194.560 ;
        RECT 30.435 194.500 30.725 194.545 ;
        RECT 22.230 194.360 30.725 194.500 ;
        RECT 13.860 194.300 14.180 194.360 ;
        RECT 19.380 194.300 19.700 194.360 ;
        RECT 28.580 194.300 28.900 194.360 ;
        RECT 30.435 194.315 30.725 194.360 ;
        RECT 33.195 194.500 33.485 194.545 ;
        RECT 33.640 194.500 33.960 194.560 ;
        RECT 33.195 194.360 33.960 194.500 ;
        RECT 33.195 194.315 33.485 194.360 ;
        RECT 33.640 194.300 33.960 194.360 ;
        RECT 37.780 194.300 38.100 194.560 ;
        RECT 38.700 194.500 39.020 194.560 ;
        RECT 41.460 194.500 41.780 194.560 ;
        RECT 38.700 194.360 41.780 194.500 ;
        RECT 38.700 194.300 39.020 194.360 ;
        RECT 41.460 194.300 41.780 194.360 ;
        RECT 8.270 193.680 43.230 194.160 ;
        RECT 8.800 193.480 9.120 193.540 ;
        RECT 23.060 193.480 23.380 193.540 ;
        RECT 24.915 193.480 25.205 193.525 ;
        RECT 8.800 193.340 20.070 193.480 ;
        RECT 8.800 193.280 9.120 193.340 ;
        RECT 9.260 193.140 9.580 193.200 ;
        RECT 17.080 193.140 17.400 193.200 ;
        RECT 9.260 193.000 17.400 193.140 ;
        RECT 9.260 192.940 9.580 193.000 ;
        RECT 10.640 192.800 10.960 192.860 ;
        RECT 10.640 192.660 14.090 192.800 ;
        RECT 10.640 192.600 10.960 192.660 ;
        RECT 11.100 192.260 11.420 192.520 ;
        RECT 12.940 192.260 13.260 192.520 ;
        RECT 13.950 192.505 14.090 192.660 ;
        RECT 14.870 192.505 15.010 193.000 ;
        RECT 17.080 192.940 17.400 193.000 ;
        RECT 15.700 192.800 16.020 192.860 ;
        RECT 15.700 192.660 19.150 192.800 ;
        RECT 15.700 192.600 16.020 192.660 ;
        RECT 13.875 192.275 14.165 192.505 ;
        RECT 14.795 192.275 15.085 192.505 ;
        RECT 16.175 192.340 16.465 192.385 ;
        RECT 9.260 192.120 9.580 192.180 ;
        RECT 11.190 192.120 11.330 192.260 ;
        RECT 16.175 192.200 16.850 192.340 ;
        RECT 18.000 192.260 18.320 192.520 ;
        RECT 18.460 192.260 18.780 192.520 ;
        RECT 19.010 192.505 19.150 192.660 ;
        RECT 19.930 192.505 20.070 193.340 ;
        RECT 23.060 193.340 25.205 193.480 ;
        RECT 23.060 193.280 23.380 193.340 ;
        RECT 24.915 193.295 25.205 193.340 ;
        RECT 27.660 193.480 27.980 193.540 ;
        RECT 29.515 193.480 29.805 193.525 ;
        RECT 35.020 193.480 35.340 193.540 ;
        RECT 27.660 193.340 29.805 193.480 ;
        RECT 27.660 193.280 27.980 193.340 ;
        RECT 29.515 193.295 29.805 193.340 ;
        RECT 31.430 193.340 35.340 193.480 ;
        RECT 31.430 193.140 31.570 193.340 ;
        RECT 35.020 193.280 35.340 193.340 ;
        RECT 41.015 193.480 41.305 193.525 ;
        RECT 43.300 193.480 43.620 193.540 ;
        RECT 41.015 193.340 43.620 193.480 ;
        RECT 41.015 193.295 41.305 193.340 ;
        RECT 43.300 193.280 43.620 193.340 ;
        RECT 22.230 193.000 31.570 193.140 ;
        RECT 31.765 193.140 32.055 193.185 ;
        RECT 33.655 193.140 33.945 193.185 ;
        RECT 36.775 193.140 37.065 193.185 ;
        RECT 31.765 193.000 37.065 193.140 ;
        RECT 22.230 192.505 22.370 193.000 ;
        RECT 31.765 192.955 32.055 193.000 ;
        RECT 33.655 192.955 33.945 193.000 ;
        RECT 36.775 192.955 37.065 193.000 ;
        RECT 39.620 193.140 39.940 193.200 ;
        RECT 41.460 193.140 41.780 193.200 ;
        RECT 39.620 193.000 41.780 193.140 ;
        RECT 39.620 192.940 39.940 193.000 ;
        RECT 41.460 192.940 41.780 193.000 ;
        RECT 30.895 192.800 31.185 192.845 ;
        RECT 35.940 192.800 36.260 192.860 ;
        RECT 30.895 192.660 36.260 192.800 ;
        RECT 30.895 192.615 31.185 192.660 ;
        RECT 35.940 192.600 36.260 192.660 ;
        RECT 18.935 192.275 19.225 192.505 ;
        RECT 19.855 192.460 20.145 192.505 ;
        RECT 22.155 192.460 22.445 192.505 ;
        RECT 19.855 192.320 22.445 192.460 ;
        RECT 19.855 192.275 20.145 192.320 ;
        RECT 22.155 192.275 22.445 192.320 ;
        RECT 22.600 192.460 22.920 192.520 ;
        RECT 27.675 192.460 27.965 192.505 ;
        RECT 28.595 192.460 28.885 192.505 ;
        RECT 22.600 192.320 28.885 192.460 ;
        RECT 22.600 192.260 22.920 192.320 ;
        RECT 27.675 192.275 27.965 192.320 ;
        RECT 28.595 192.275 28.885 192.320 ;
        RECT 31.360 192.460 31.650 192.505 ;
        RECT 33.195 192.460 33.485 192.505 ;
        RECT 36.775 192.460 37.065 192.505 ;
        RECT 31.360 192.320 37.065 192.460 ;
        RECT 31.360 192.275 31.650 192.320 ;
        RECT 33.195 192.275 33.485 192.320 ;
        RECT 36.775 192.275 37.065 192.320 ;
        RECT 13.415 192.120 13.705 192.165 ;
        RECT 16.175 192.155 16.465 192.200 ;
        RECT 16.710 192.120 16.850 192.200 ;
        RECT 23.520 192.120 23.840 192.180 ;
        RECT 23.995 192.120 24.285 192.165 ;
        RECT 9.260 191.980 13.705 192.120 ;
        RECT 9.260 191.920 9.580 191.980 ;
        RECT 13.415 191.935 13.705 191.980 ;
        RECT 13.950 191.980 15.930 192.120 ;
        RECT 16.710 191.980 18.690 192.120 ;
        RECT 11.100 191.780 11.420 191.840 ;
        RECT 12.035 191.780 12.325 191.825 ;
        RECT 11.100 191.640 12.325 191.780 ;
        RECT 11.100 191.580 11.420 191.640 ;
        RECT 12.035 191.595 12.325 191.640 ;
        RECT 12.940 191.780 13.260 191.840 ;
        RECT 13.950 191.780 14.090 191.980 ;
        RECT 12.940 191.640 14.090 191.780 ;
        RECT 14.780 191.780 15.100 191.840 ;
        RECT 15.255 191.780 15.545 191.825 ;
        RECT 14.780 191.640 15.545 191.780 ;
        RECT 15.790 191.780 15.930 191.980 ;
        RECT 17.095 191.780 17.385 191.825 ;
        RECT 15.790 191.640 17.385 191.780 ;
        RECT 18.550 191.780 18.690 191.980 ;
        RECT 23.520 191.980 24.285 192.120 ;
        RECT 23.520 191.920 23.840 191.980 ;
        RECT 23.995 191.935 24.285 191.980 ;
        RECT 26.280 191.920 26.600 192.180 ;
        RECT 32.260 191.920 32.580 192.180 ;
        RECT 37.855 192.165 38.145 192.480 ;
        RECT 40.095 192.460 40.385 192.505 ;
        RECT 41.920 192.460 42.240 192.520 ;
        RECT 40.095 192.320 42.240 192.460 ;
        RECT 40.095 192.275 40.385 192.320 ;
        RECT 41.920 192.260 42.240 192.320 ;
        RECT 34.555 192.120 35.205 192.165 ;
        RECT 37.855 192.120 38.445 192.165 ;
        RECT 32.810 191.980 38.445 192.120 ;
        RECT 18.920 191.780 19.240 191.840 ;
        RECT 18.550 191.640 19.240 191.780 ;
        RECT 26.370 191.780 26.510 191.920 ;
        RECT 28.580 191.780 28.900 191.840 ;
        RECT 32.810 191.780 32.950 191.980 ;
        RECT 34.555 191.935 35.205 191.980 ;
        RECT 38.155 191.935 38.445 191.980 ;
        RECT 26.370 191.640 32.950 191.780 ;
        RECT 33.640 191.780 33.960 191.840 ;
        RECT 35.940 191.780 36.260 191.840 ;
        RECT 33.640 191.640 36.260 191.780 ;
        RECT 12.940 191.580 13.260 191.640 ;
        RECT 14.780 191.580 15.100 191.640 ;
        RECT 15.255 191.595 15.545 191.640 ;
        RECT 17.095 191.595 17.385 191.640 ;
        RECT 18.920 191.580 19.240 191.640 ;
        RECT 28.580 191.580 28.900 191.640 ;
        RECT 33.640 191.580 33.960 191.640 ;
        RECT 35.940 191.580 36.260 191.640 ;
        RECT 36.860 191.780 37.180 191.840 ;
        RECT 39.635 191.780 39.925 191.825 ;
        RECT 36.860 191.640 39.925 191.780 ;
        RECT 36.860 191.580 37.180 191.640 ;
        RECT 39.635 191.595 39.925 191.640 ;
        RECT 8.270 190.960 43.230 191.440 ;
        RECT 13.860 190.760 14.180 190.820 ;
        RECT 13.860 190.620 15.930 190.760 ;
        RECT 13.860 190.560 14.180 190.620 ;
        RECT 11.575 190.420 11.865 190.465 ;
        RECT 12.940 190.420 13.260 190.480 ;
        RECT 15.790 190.465 15.930 190.620 ;
        RECT 22.600 190.560 22.920 190.820 ;
        RECT 34.560 190.760 34.880 190.820 ;
        RECT 35.035 190.760 35.325 190.805 ;
        RECT 34.560 190.620 35.325 190.760 ;
        RECT 34.560 190.560 34.880 190.620 ;
        RECT 35.035 190.575 35.325 190.620 ;
        RECT 36.875 190.760 37.165 190.805 ;
        RECT 40.080 190.760 40.400 190.820 ;
        RECT 36.875 190.620 40.400 190.760 ;
        RECT 36.875 190.575 37.165 190.620 ;
        RECT 40.080 190.560 40.400 190.620 ;
        RECT 11.575 190.280 13.260 190.420 ;
        RECT 11.575 190.235 11.865 190.280 ;
        RECT 12.940 190.220 13.260 190.280 ;
        RECT 15.715 190.235 16.005 190.465 ;
        RECT 10.640 190.080 10.960 190.140 ;
        RECT 12.495 190.080 12.785 190.125 ;
        RECT 10.640 189.940 12.785 190.080 ;
        RECT 10.640 189.880 10.960 189.940 ;
        RECT 12.495 189.895 12.785 189.940 ;
        RECT 14.675 190.080 14.965 190.125 ;
        RECT 14.675 189.895 15.010 190.080 ;
        RECT 9.260 189.540 9.580 189.800 ;
        RECT 14.870 189.740 15.010 189.895 ;
        RECT 15.240 189.880 15.560 190.140 ;
        RECT 16.620 189.880 16.940 190.140 ;
        RECT 17.555 190.080 17.845 190.125 ;
        RECT 19.380 190.080 19.700 190.140 ;
        RECT 17.555 189.940 19.700 190.080 ;
        RECT 17.555 189.895 17.845 189.940 ;
        RECT 19.380 189.880 19.700 189.940 ;
        RECT 22.155 189.895 22.445 190.125 ;
        RECT 22.690 190.080 22.830 190.560 ;
        RECT 33.655 190.420 33.945 190.465 ;
        RECT 41.000 190.420 41.320 190.480 ;
        RECT 33.655 190.280 41.320 190.420 ;
        RECT 33.655 190.235 33.945 190.280 ;
        RECT 41.000 190.220 41.320 190.280 ;
        RECT 22.690 189.940 23.290 190.080 ;
        RECT 18.000 189.740 18.320 189.800 ;
        RECT 14.870 189.600 18.320 189.740 ;
        RECT 18.000 189.540 18.320 189.600 ;
        RECT 9.350 189.400 9.490 189.540 ;
        RECT 15.240 189.400 15.560 189.460 ;
        RECT 9.350 189.260 15.560 189.400 ;
        RECT 15.240 189.200 15.560 189.260 ;
        RECT 18.460 189.200 18.780 189.460 ;
        RECT 7.420 189.060 7.740 189.120 ;
        RECT 10.195 189.060 10.485 189.105 ;
        RECT 7.420 188.920 10.485 189.060 ;
        RECT 7.420 188.860 7.740 188.920 ;
        RECT 10.195 188.875 10.485 188.920 ;
        RECT 13.400 188.860 13.720 189.120 ;
        RECT 13.860 188.860 14.180 189.120 ;
        RECT 18.000 189.060 18.320 189.120 ;
        RECT 20.315 189.060 20.605 189.105 ;
        RECT 18.000 188.920 20.605 189.060 ;
        RECT 22.230 189.060 22.370 189.895 ;
        RECT 23.150 189.785 23.290 189.940 ;
        RECT 35.955 189.895 36.245 190.125 ;
        RECT 22.615 189.555 22.905 189.785 ;
        RECT 23.075 189.555 23.365 189.785 ;
        RECT 22.690 189.400 22.830 189.555 ;
        RECT 32.260 189.400 32.580 189.460 ;
        RECT 36.030 189.400 36.170 189.895 ;
        RECT 39.620 189.880 39.940 190.140 ;
        RECT 41.475 190.080 41.765 190.125 ;
        RECT 43.300 190.080 43.620 190.140 ;
        RECT 41.475 189.940 43.620 190.080 ;
        RECT 41.475 189.895 41.765 189.940 ;
        RECT 43.300 189.880 43.620 189.940 ;
        RECT 60.960 189.895 61.340 190.245 ;
        RECT 22.690 189.260 36.170 189.400 ;
        RECT 32.260 189.200 32.580 189.260 ;
        RECT 23.520 189.060 23.840 189.120 ;
        RECT 22.230 188.920 23.840 189.060 ;
        RECT 18.000 188.860 18.320 188.920 ;
        RECT 20.315 188.875 20.605 188.920 ;
        RECT 23.520 188.860 23.840 188.920 ;
        RECT 25.820 189.060 26.140 189.120 ;
        RECT 26.295 189.060 26.585 189.105 ;
        RECT 25.820 188.920 26.585 189.060 ;
        RECT 25.820 188.860 26.140 188.920 ;
        RECT 26.295 188.875 26.585 188.920 ;
        RECT 31.800 189.060 32.120 189.120 ;
        RECT 40.555 189.060 40.845 189.105 ;
        RECT 41.000 189.060 41.320 189.120 ;
        RECT 31.800 188.920 41.320 189.060 ;
        RECT 31.800 188.860 32.120 188.920 ;
        RECT 40.555 188.875 40.845 188.920 ;
        RECT 41.000 188.860 41.320 188.920 ;
        RECT 8.270 188.240 43.230 188.720 ;
        RECT 58.510 188.210 59.890 188.285 ;
        RECT 18.000 187.840 18.320 188.100 ;
        RECT 25.375 188.040 25.665 188.085 ;
        RECT 27.200 188.040 27.520 188.100 ;
        RECT 25.375 187.900 27.520 188.040 ;
        RECT 25.375 187.855 25.665 187.900 ;
        RECT 27.200 187.840 27.520 187.900 ;
        RECT 36.400 187.840 36.720 188.100 ;
        RECT 55.245 187.860 59.890 188.210 ;
        RECT 15.715 187.700 16.005 187.745 ;
        RECT 17.080 187.700 17.400 187.760 ;
        RECT 18.090 187.700 18.230 187.840 ;
        RECT 23.520 187.700 23.840 187.760 ;
        RECT 15.715 187.560 17.400 187.700 ;
        RECT 15.715 187.515 16.005 187.560 ;
        RECT 17.080 187.500 17.400 187.560 ;
        RECT 17.630 187.560 18.230 187.700 ;
        RECT 22.230 187.560 23.840 187.700 ;
        RECT 13.860 187.160 14.180 187.420 ;
        RECT 11.100 187.020 11.420 187.080 ;
        RECT 11.575 187.020 11.865 187.065 ;
        RECT 11.100 186.880 11.865 187.020 ;
        RECT 13.950 187.020 14.090 187.160 ;
        RECT 14.335 187.020 14.625 187.065 ;
        RECT 13.950 186.880 14.625 187.020 ;
        RECT 11.100 186.820 11.420 186.880 ;
        RECT 11.575 186.835 11.865 186.880 ;
        RECT 14.335 186.835 14.625 186.880 ;
        RECT 16.635 187.020 16.925 187.065 ;
        RECT 17.630 187.020 17.770 187.560 ;
        RECT 19.855 187.360 20.145 187.405 ;
        RECT 16.635 186.880 17.770 187.020 ;
        RECT 18.090 187.220 20.145 187.360 ;
        RECT 16.635 186.835 16.925 186.880 ;
        RECT 9.720 186.480 10.040 186.740 ;
        RECT 12.480 186.480 12.800 186.740 ;
        RECT 12.940 186.680 13.260 186.740 ;
        RECT 18.090 186.680 18.230 187.220 ;
        RECT 19.855 187.175 20.145 187.220 ;
        RECT 18.920 186.820 19.240 187.080 ;
        RECT 19.010 186.680 19.150 186.820 ;
        RECT 12.940 186.540 18.230 186.680 ;
        RECT 18.550 186.540 19.150 186.680 ;
        RECT 12.940 186.480 13.260 186.540 ;
        RECT 17.095 186.340 17.385 186.385 ;
        RECT 18.550 186.340 18.690 186.540 ;
        RECT 22.230 186.400 22.370 187.560 ;
        RECT 23.520 187.500 23.840 187.560 ;
        RECT 22.600 187.160 22.920 187.420 ;
        RECT 34.560 187.360 34.880 187.420 ;
        RECT 23.610 187.220 34.880 187.360 ;
        RECT 23.610 187.065 23.750 187.220 ;
        RECT 34.560 187.160 34.880 187.220 ;
        RECT 36.860 187.360 37.180 187.420 ;
        RECT 40.080 187.360 40.400 187.420 ;
        RECT 41.015 187.360 41.305 187.405 ;
        RECT 36.860 187.220 41.305 187.360 ;
        RECT 36.860 187.160 37.180 187.220 ;
        RECT 40.080 187.160 40.400 187.220 ;
        RECT 41.015 187.175 41.305 187.220 ;
        RECT 23.535 186.835 23.825 187.065 ;
        RECT 25.360 186.820 25.680 187.080 ;
        RECT 29.055 187.020 29.345 187.065 ;
        RECT 25.910 186.880 29.345 187.020 ;
        RECT 23.075 186.680 23.365 186.725 ;
        RECT 25.450 186.680 25.590 186.820 ;
        RECT 25.910 186.740 26.050 186.880 ;
        RECT 29.055 186.835 29.345 186.880 ;
        RECT 23.075 186.540 25.590 186.680 ;
        RECT 23.075 186.495 23.365 186.540 ;
        RECT 25.820 186.480 26.140 186.740 ;
        RECT 26.755 186.495 27.045 186.725 ;
        RECT 28.595 186.680 28.885 186.725 ;
        RECT 44.680 186.680 45.000 186.740 ;
        RECT 28.595 186.540 45.000 186.680 ;
        RECT 28.595 186.495 28.885 186.540 ;
        RECT 17.095 186.200 18.690 186.340 ;
        RECT 17.095 186.155 17.385 186.200 ;
        RECT 18.920 186.140 19.240 186.400 ;
        RECT 19.395 186.340 19.685 186.385 ;
        RECT 22.140 186.340 22.460 186.400 ;
        RECT 19.395 186.200 22.460 186.340 ;
        RECT 19.395 186.155 19.685 186.200 ;
        RECT 22.140 186.140 22.460 186.200 ;
        RECT 23.520 186.340 23.840 186.400 ;
        RECT 26.830 186.340 26.970 186.495 ;
        RECT 44.680 186.480 45.000 186.540 ;
        RECT 23.520 186.200 26.970 186.340 ;
        RECT 31.800 186.340 32.120 186.400 ;
        RECT 38.255 186.340 38.545 186.385 ;
        RECT 31.800 186.200 38.545 186.340 ;
        RECT 23.520 186.140 23.840 186.200 ;
        RECT 31.800 186.140 32.120 186.200 ;
        RECT 38.255 186.155 38.545 186.200 ;
        RECT 8.270 185.520 43.230 186.000 ;
        RECT 9.260 185.120 9.580 185.380 ;
        RECT 10.640 185.320 10.960 185.380 ;
        RECT 19.840 185.320 20.160 185.380 ;
        RECT 30.880 185.320 31.200 185.380 ;
        RECT 10.640 185.180 20.160 185.320 ;
        RECT 10.640 185.120 10.960 185.180 ;
        RECT 19.840 185.120 20.160 185.180 ;
        RECT 25.910 185.180 31.200 185.320 ;
        RECT 9.350 184.980 9.490 185.120 ;
        RECT 15.720 184.980 16.010 185.025 ;
        RECT 17.580 184.980 17.870 185.025 ;
        RECT 9.350 184.840 13.630 184.980 ;
        RECT 8.800 184.640 9.120 184.700 ;
        RECT 12.035 184.640 12.325 184.685 ;
        RECT 8.800 184.500 12.325 184.640 ;
        RECT 8.800 184.440 9.120 184.500 ;
        RECT 10.730 184.360 10.870 184.500 ;
        RECT 12.035 184.455 12.325 184.500 ;
        RECT 12.495 184.640 12.785 184.685 ;
        RECT 12.940 184.640 13.260 184.700 ;
        RECT 13.490 184.685 13.630 184.840 ;
        RECT 15.720 184.840 17.870 184.980 ;
        RECT 15.720 184.795 16.010 184.840 ;
        RECT 17.580 184.795 17.870 184.840 ;
        RECT 18.500 184.980 18.790 185.025 ;
        RECT 21.760 184.980 22.050 185.025 ;
        RECT 23.980 184.980 24.300 185.040 ;
        RECT 25.910 185.025 26.050 185.180 ;
        RECT 30.880 185.120 31.200 185.180 ;
        RECT 32.260 185.320 32.580 185.380 ;
        RECT 33.195 185.320 33.485 185.365 ;
        RECT 32.260 185.180 33.485 185.320 ;
        RECT 32.260 185.120 32.580 185.180 ;
        RECT 33.195 185.135 33.485 185.180 ;
        RECT 28.580 185.025 28.900 185.040 ;
        RECT 18.500 184.840 24.300 184.980 ;
        RECT 18.500 184.795 18.790 184.840 ;
        RECT 21.760 184.795 22.050 184.840 ;
        RECT 12.495 184.500 13.260 184.640 ;
        RECT 12.495 184.455 12.785 184.500 ;
        RECT 10.640 184.100 10.960 184.360 ;
        RECT 11.100 184.300 11.420 184.360 ;
        RECT 12.570 184.300 12.710 184.455 ;
        RECT 12.940 184.440 13.260 184.500 ;
        RECT 13.415 184.455 13.705 184.685 ;
        RECT 17.655 184.640 17.870 184.795 ;
        RECT 23.980 184.780 24.300 184.840 ;
        RECT 25.835 184.795 26.125 185.025 ;
        RECT 28.115 184.980 28.900 185.025 ;
        RECT 31.715 184.980 32.005 185.025 ;
        RECT 28.115 184.840 32.005 184.980 ;
        RECT 28.115 184.795 28.900 184.840 ;
        RECT 28.580 184.780 28.900 184.795 ;
        RECT 31.415 184.795 32.005 184.840 ;
        RECT 19.900 184.640 20.190 184.685 ;
        RECT 14.870 184.500 17.310 184.640 ;
        RECT 17.655 184.500 20.190 184.640 ;
        RECT 11.100 184.160 12.710 184.300 ;
        RECT 13.860 184.300 14.180 184.360 ;
        RECT 14.870 184.345 15.010 184.500 ;
        RECT 14.795 184.300 15.085 184.345 ;
        RECT 13.860 184.160 15.085 184.300 ;
        RECT 11.100 184.100 11.420 184.160 ;
        RECT 13.860 184.100 14.180 184.160 ;
        RECT 14.795 184.115 15.085 184.160 ;
        RECT 16.620 184.100 16.940 184.360 ;
        RECT 17.170 184.300 17.310 184.500 ;
        RECT 19.900 184.455 20.190 184.500 ;
        RECT 24.455 184.455 24.745 184.685 ;
        RECT 24.920 184.640 25.210 184.685 ;
        RECT 26.755 184.640 27.045 184.685 ;
        RECT 30.335 184.640 30.625 184.685 ;
        RECT 24.920 184.500 30.625 184.640 ;
        RECT 24.920 184.455 25.210 184.500 ;
        RECT 26.755 184.455 27.045 184.500 ;
        RECT 30.335 184.455 30.625 184.500 ;
        RECT 31.415 184.480 31.705 184.795 ;
        RECT 33.270 184.640 33.410 185.135 ;
        RECT 34.560 185.120 34.880 185.380 ;
        RECT 40.080 185.120 40.400 185.380 ;
        RECT 40.540 185.320 40.860 185.380 ;
        RECT 41.475 185.320 41.765 185.365 ;
        RECT 40.540 185.180 41.765 185.320 ;
        RECT 40.540 185.120 40.860 185.180 ;
        RECT 41.475 185.135 41.765 185.180 ;
        RECT 39.620 184.780 39.940 185.040 ;
        RECT 40.170 184.980 40.310 185.120 ;
        RECT 40.170 184.840 40.770 184.980 ;
        RECT 40.630 184.685 40.770 184.840 ;
        RECT 43.760 184.780 44.080 185.040 ;
        RECT 37.335 184.640 37.625 184.685 ;
        RECT 33.270 184.500 37.625 184.640 ;
        RECT 37.335 184.455 37.625 184.500 ;
        RECT 38.715 184.455 39.005 184.685 ;
        RECT 40.095 184.455 40.385 184.685 ;
        RECT 40.555 184.640 40.845 184.685 ;
        RECT 41.460 184.640 41.780 184.700 ;
        RECT 40.555 184.500 41.780 184.640 ;
        RECT 40.555 184.455 40.845 184.500 ;
        RECT 17.540 184.300 17.860 184.360 ;
        RECT 24.530 184.300 24.670 184.455 ;
        RECT 17.170 184.160 24.670 184.300 ;
        RECT 35.020 184.300 35.340 184.360 ;
        RECT 36.860 184.300 37.180 184.360 ;
        RECT 38.790 184.300 38.930 184.455 ;
        RECT 35.020 184.160 38.930 184.300 ;
        RECT 40.170 184.300 40.310 184.455 ;
        RECT 41.460 184.440 41.780 184.500 ;
        RECT 41.920 184.300 42.240 184.360 ;
        RECT 43.850 184.300 43.990 184.780 ;
        RECT 40.170 184.160 43.990 184.300 ;
        RECT 17.540 184.100 17.860 184.160 ;
        RECT 35.020 184.100 35.340 184.160 ;
        RECT 36.860 184.100 37.180 184.160 ;
        RECT 41.920 184.100 42.240 184.160 ;
        RECT 15.260 183.960 15.550 184.005 ;
        RECT 17.120 183.960 17.410 184.005 ;
        RECT 19.900 183.960 20.190 184.005 ;
        RECT 15.260 183.820 20.190 183.960 ;
        RECT 15.260 183.775 15.550 183.820 ;
        RECT 17.120 183.775 17.410 183.820 ;
        RECT 19.900 183.775 20.190 183.820 ;
        RECT 25.325 183.960 25.615 184.005 ;
        RECT 27.215 183.960 27.505 184.005 ;
        RECT 30.335 183.960 30.625 184.005 ;
        RECT 25.325 183.820 30.625 183.960 ;
        RECT 25.325 183.775 25.615 183.820 ;
        RECT 27.215 183.775 27.505 183.820 ;
        RECT 30.335 183.775 30.625 183.820 ;
        RECT 2.820 183.620 3.140 183.680 ;
        RECT 12.480 183.620 12.800 183.680 ;
        RECT 2.820 183.480 12.800 183.620 ;
        RECT 2.820 183.420 3.140 183.480 ;
        RECT 12.480 183.420 12.800 183.480 ;
        RECT 14.335 183.620 14.625 183.665 ;
        RECT 19.380 183.620 19.700 183.680 ;
        RECT 14.335 183.480 19.700 183.620 ;
        RECT 14.335 183.435 14.625 183.480 ;
        RECT 19.380 183.420 19.700 183.480 ;
        RECT 22.140 183.620 22.460 183.680 ;
        RECT 23.765 183.620 24.055 183.665 ;
        RECT 28.120 183.620 28.440 183.680 ;
        RECT 22.140 183.480 28.440 183.620 ;
        RECT 22.140 183.420 22.460 183.480 ;
        RECT 23.765 183.435 24.055 183.480 ;
        RECT 28.120 183.420 28.440 183.480 ;
        RECT 35.020 183.620 35.340 183.680 ;
        RECT 41.000 183.620 41.320 183.680 ;
        RECT 35.020 183.480 41.320 183.620 ;
        RECT 35.020 183.420 35.340 183.480 ;
        RECT 41.000 183.420 41.320 183.480 ;
        RECT 8.270 182.800 43.230 183.280 ;
        RECT 10.180 182.600 10.500 182.660 ;
        RECT 34.560 182.600 34.880 182.660 ;
        RECT 10.180 182.460 34.880 182.600 ;
        RECT 10.180 182.400 10.500 182.460 ;
        RECT 34.560 182.400 34.880 182.460 ;
        RECT 40.540 182.600 40.860 182.660 ;
        RECT 41.015 182.600 41.305 182.645 ;
        RECT 40.540 182.460 41.305 182.600 ;
        RECT 40.540 182.400 40.860 182.460 ;
        RECT 41.015 182.415 41.305 182.460 ;
        RECT 12.905 182.260 13.195 182.305 ;
        RECT 14.795 182.260 15.085 182.305 ;
        RECT 17.915 182.260 18.205 182.305 ;
        RECT 12.905 182.120 18.205 182.260 ;
        RECT 12.905 182.075 13.195 182.120 ;
        RECT 14.795 182.075 15.085 182.120 ;
        RECT 17.915 182.075 18.205 182.120 ;
        RECT 25.935 182.260 26.225 182.305 ;
        RECT 29.055 182.260 29.345 182.305 ;
        RECT 30.945 182.260 31.235 182.305 ;
        RECT 25.935 182.120 31.235 182.260 ;
        RECT 25.935 182.075 26.225 182.120 ;
        RECT 29.055 182.075 29.345 182.120 ;
        RECT 30.945 182.075 31.235 182.120 ;
        RECT 33.145 182.260 33.435 182.305 ;
        RECT 35.035 182.260 35.325 182.305 ;
        RECT 38.155 182.260 38.445 182.305 ;
        RECT 33.145 182.120 38.445 182.260 ;
        RECT 33.145 182.075 33.435 182.120 ;
        RECT 35.035 182.075 35.325 182.120 ;
        RECT 38.155 182.075 38.445 182.120 ;
        RECT 12.035 181.920 12.325 181.965 ;
        RECT 13.860 181.920 14.180 181.980 ;
        RECT 12.035 181.780 14.180 181.920 ;
        RECT 12.035 181.735 12.325 181.780 ;
        RECT 13.860 181.720 14.180 181.780 ;
        RECT 17.080 181.920 17.400 181.980 ;
        RECT 23.980 181.920 24.300 181.980 ;
        RECT 28.580 181.920 28.900 181.980 ;
        RECT 17.080 181.780 28.900 181.920 ;
        RECT 17.080 181.720 17.400 181.780 ;
        RECT 12.500 181.580 12.790 181.625 ;
        RECT 14.335 181.580 14.625 181.625 ;
        RECT 17.915 181.580 18.205 181.625 ;
        RECT 19.010 181.600 19.150 181.780 ;
        RECT 23.980 181.720 24.300 181.780 ;
        RECT 12.500 181.440 18.205 181.580 ;
        RECT 12.500 181.395 12.790 181.440 ;
        RECT 14.335 181.395 14.625 181.440 ;
        RECT 17.915 181.395 18.205 181.440 ;
        RECT 13.415 181.240 13.705 181.285 ;
        RECT 14.780 181.240 15.100 181.300 ;
        RECT 18.995 181.285 19.285 181.600 ;
        RECT 21.680 181.380 22.000 181.640 ;
        RECT 23.060 181.380 23.380 181.640 ;
        RECT 24.990 181.600 25.130 181.780 ;
        RECT 28.580 181.720 28.900 181.780 ;
        RECT 31.815 181.920 32.105 181.965 ;
        RECT 32.275 181.920 32.565 181.965 ;
        RECT 36.400 181.920 36.720 181.980 ;
        RECT 31.815 181.780 36.720 181.920 ;
        RECT 31.815 181.735 32.105 181.780 ;
        RECT 32.275 181.735 32.565 181.780 ;
        RECT 36.400 181.720 36.720 181.780 ;
        RECT 13.415 181.100 15.100 181.240 ;
        RECT 13.415 181.055 13.705 181.100 ;
        RECT 14.780 181.040 15.100 181.100 ;
        RECT 15.695 181.240 16.345 181.285 ;
        RECT 18.995 181.240 19.585 181.285 ;
        RECT 23.150 181.240 23.290 181.380 ;
        RECT 24.855 181.285 25.145 181.600 ;
        RECT 25.935 181.580 26.225 181.625 ;
        RECT 29.515 181.580 29.805 181.625 ;
        RECT 31.350 181.580 31.640 181.625 ;
        RECT 25.935 181.440 31.640 181.580 ;
        RECT 25.935 181.395 26.225 181.440 ;
        RECT 29.515 181.395 29.805 181.440 ;
        RECT 31.350 181.395 31.640 181.440 ;
        RECT 32.740 181.580 33.030 181.625 ;
        RECT 34.575 181.580 34.865 181.625 ;
        RECT 38.155 181.580 38.445 181.625 ;
        RECT 32.740 181.440 38.445 181.580 ;
        RECT 32.740 181.395 33.030 181.440 ;
        RECT 34.575 181.395 34.865 181.440 ;
        RECT 38.155 181.395 38.445 181.440 ;
        RECT 15.695 181.100 19.585 181.240 ;
        RECT 15.695 181.055 16.345 181.100 ;
        RECT 19.295 181.055 19.585 181.100 ;
        RECT 20.850 181.100 23.290 181.240 ;
        RECT 24.555 181.240 25.145 181.285 ;
        RECT 27.795 181.240 28.445 181.285 ;
        RECT 24.555 181.100 28.445 181.240 ;
        RECT 20.850 180.960 20.990 181.100 ;
        RECT 24.555 181.055 24.845 181.100 ;
        RECT 27.795 181.055 28.445 181.100 ;
        RECT 30.435 181.240 30.725 181.285 ;
        RECT 31.800 181.240 32.120 181.300 ;
        RECT 30.435 181.100 32.120 181.240 ;
        RECT 30.435 181.055 30.725 181.100 ;
        RECT 31.800 181.040 32.120 181.100 ;
        RECT 32.260 181.240 32.580 181.300 ;
        RECT 33.655 181.240 33.945 181.285 ;
        RECT 32.260 181.100 33.945 181.240 ;
        RECT 32.260 181.040 32.580 181.100 ;
        RECT 33.655 181.055 33.945 181.100 ;
        RECT 35.020 181.240 35.340 181.300 ;
        RECT 39.235 181.285 39.525 181.600 ;
        RECT 35.935 181.240 36.585 181.285 ;
        RECT 39.235 181.240 39.825 181.285 ;
        RECT 35.020 181.100 39.825 181.240 ;
        RECT 35.020 181.040 35.340 181.100 ;
        RECT 35.935 181.055 36.585 181.100 ;
        RECT 39.535 181.055 39.825 181.100 ;
        RECT 40.080 181.240 40.400 181.300 ;
        RECT 41.460 181.240 41.780 181.300 ;
        RECT 40.080 181.100 41.780 181.240 ;
        RECT 40.080 181.040 40.400 181.100 ;
        RECT 41.460 181.040 41.780 181.100 ;
        RECT 41.920 181.040 42.240 181.300 ;
        RECT 18.460 180.900 18.780 180.960 ;
        RECT 20.760 180.900 21.080 180.960 ;
        RECT 18.460 180.760 21.080 180.900 ;
        RECT 18.460 180.700 18.780 180.760 ;
        RECT 20.760 180.700 21.080 180.760 ;
        RECT 22.600 180.700 22.920 180.960 ;
        RECT 23.075 180.900 23.365 180.945 ;
        RECT 29.040 180.900 29.360 180.960 ;
        RECT 23.075 180.760 29.360 180.900 ;
        RECT 23.075 180.715 23.365 180.760 ;
        RECT 29.040 180.700 29.360 180.760 ;
        RECT 38.240 180.900 38.560 180.960 ;
        RECT 42.010 180.900 42.150 181.040 ;
        RECT 38.240 180.760 42.150 180.900 ;
        RECT 38.240 180.700 38.560 180.760 ;
        RECT 8.270 180.080 43.230 180.560 ;
        RECT 11.100 179.880 11.420 179.940 ;
        RECT 13.415 179.880 13.705 179.925 ;
        RECT 14.780 179.880 15.100 179.940 ;
        RECT 11.100 179.740 15.100 179.880 ;
        RECT 11.100 179.680 11.420 179.740 ;
        RECT 13.415 179.695 13.705 179.740 ;
        RECT 14.780 179.680 15.100 179.740 ;
        RECT 15.255 179.880 15.545 179.925 ;
        RECT 19.840 179.880 20.160 179.940 ;
        RECT 24.915 179.880 25.205 179.925 ;
        RECT 15.255 179.740 19.610 179.880 ;
        RECT 15.255 179.695 15.545 179.740 ;
        RECT 19.470 179.540 19.610 179.740 ;
        RECT 19.840 179.740 25.205 179.880 ;
        RECT 19.840 179.680 20.160 179.740 ;
        RECT 24.915 179.695 25.205 179.740 ;
        RECT 26.280 179.880 26.600 179.940 ;
        RECT 26.755 179.880 27.045 179.925 ;
        RECT 26.280 179.740 27.045 179.880 ;
        RECT 26.280 179.680 26.600 179.740 ;
        RECT 26.755 179.695 27.045 179.740 ;
        RECT 32.260 179.680 32.580 179.940 ;
        RECT 34.560 179.880 34.880 179.940 ;
        RECT 38.255 179.880 38.545 179.925 ;
        RECT 34.560 179.740 38.545 179.880 ;
        RECT 34.560 179.680 34.880 179.740 ;
        RECT 38.255 179.695 38.545 179.740 ;
        RECT 40.080 179.680 40.400 179.940 ;
        RECT 23.520 179.540 23.840 179.600 ;
        RECT 12.110 179.400 16.390 179.540 ;
        RECT 19.470 179.400 23.840 179.540 ;
        RECT 12.110 179.245 12.250 179.400 ;
        RECT 12.035 179.015 12.325 179.245 ;
        RECT 12.940 179.000 13.260 179.260 ;
        RECT 14.335 179.200 14.625 179.245 ;
        RECT 13.490 179.060 14.625 179.200 ;
        RECT 10.640 178.860 10.960 178.920 ;
        RECT 13.490 178.860 13.630 179.060 ;
        RECT 14.335 179.015 14.625 179.060 ;
        RECT 10.640 178.720 13.630 178.860 ;
        RECT 13.860 178.860 14.180 178.920 ;
        RECT 15.715 178.860 16.005 178.905 ;
        RECT 13.860 178.720 16.005 178.860 ;
        RECT 16.250 178.860 16.390 179.400 ;
        RECT 23.520 179.340 23.840 179.400 ;
        RECT 24.455 179.540 24.745 179.585 ;
        RECT 25.820 179.540 26.140 179.600 ;
        RECT 24.455 179.400 26.140 179.540 ;
        RECT 24.455 179.355 24.745 179.400 ;
        RECT 25.820 179.340 26.140 179.400 ;
        RECT 35.480 179.340 35.800 179.600 ;
        RECT 36.860 179.540 37.180 179.600 ;
        RECT 40.170 179.540 40.310 179.680 ;
        RECT 36.860 179.400 38.930 179.540 ;
        RECT 36.860 179.340 37.180 179.400 ;
        RECT 29.040 179.200 29.360 179.260 ;
        RECT 31.340 179.200 31.660 179.260 ;
        RECT 36.415 179.200 36.705 179.245 ;
        RECT 37.795 179.200 38.085 179.245 ;
        RECT 38.240 179.200 38.560 179.260 ;
        RECT 29.040 179.060 36.705 179.200 ;
        RECT 29.040 179.000 29.360 179.060 ;
        RECT 31.340 179.000 31.660 179.060 ;
        RECT 36.415 179.015 36.705 179.060 ;
        RECT 36.950 179.060 38.560 179.200 ;
        RECT 19.840 178.860 20.160 178.920 ;
        RECT 16.250 178.720 20.160 178.860 ;
        RECT 10.640 178.660 10.960 178.720 ;
        RECT 13.860 178.660 14.180 178.720 ;
        RECT 15.715 178.675 16.005 178.720 ;
        RECT 19.840 178.660 20.160 178.720 ;
        RECT 20.760 178.860 21.080 178.920 ;
        RECT 27.215 178.860 27.505 178.905 ;
        RECT 20.760 178.720 27.505 178.860 ;
        RECT 20.760 178.660 21.080 178.720 ;
        RECT 27.215 178.675 27.505 178.720 ;
        RECT 27.660 178.660 27.980 178.920 ;
        RECT 28.580 178.860 28.900 178.920 ;
        RECT 36.950 178.860 37.090 179.060 ;
        RECT 37.795 179.015 38.085 179.060 ;
        RECT 38.240 179.000 38.560 179.060 ;
        RECT 28.580 178.720 37.090 178.860 ;
        RECT 37.335 178.860 37.625 178.905 ;
        RECT 38.790 178.860 38.930 179.400 ;
        RECT 39.250 179.400 40.310 179.540 ;
        RECT 39.250 179.245 39.390 179.400 ;
        RECT 40.540 179.340 40.860 179.600 ;
        RECT 39.175 179.015 39.465 179.245 ;
        RECT 39.635 179.015 39.925 179.245 ;
        RECT 40.095 179.200 40.385 179.245 ;
        RECT 40.630 179.200 40.770 179.340 ;
        RECT 40.095 179.060 40.770 179.200 ;
        RECT 40.095 179.015 40.385 179.060 ;
        RECT 37.335 178.720 38.930 178.860 ;
        RECT 28.580 178.660 28.900 178.720 ;
        RECT 37.335 178.675 37.625 178.720 ;
        RECT 16.160 178.520 16.480 178.580 ;
        RECT 23.980 178.520 24.300 178.580 ;
        RECT 27.750 178.520 27.890 178.660 ;
        RECT 11.650 178.380 15.930 178.520 ;
        RECT 11.650 178.225 11.790 178.380 ;
        RECT 11.575 177.995 11.865 178.225 ;
        RECT 15.790 178.180 15.930 178.380 ;
        RECT 16.160 178.380 27.890 178.520 ;
        RECT 16.160 178.320 16.480 178.380 ;
        RECT 23.980 178.320 24.300 178.380 ;
        RECT 23.520 178.180 23.840 178.240 ;
        RECT 15.790 178.040 23.840 178.180 ;
        RECT 23.520 177.980 23.840 178.040 ;
        RECT 36.860 178.180 37.180 178.240 ;
        RECT 39.710 178.180 39.850 179.015 ;
        RECT 41.000 179.000 41.320 179.260 ;
        RECT 36.860 178.040 39.850 178.180 ;
        RECT 36.860 177.980 37.180 178.040 ;
        RECT 8.270 177.360 43.230 177.840 ;
        RECT 21.695 177.160 21.985 177.205 ;
        RECT 22.600 177.160 22.920 177.220 ;
        RECT 21.695 177.020 22.920 177.160 ;
        RECT 21.695 176.975 21.985 177.020 ;
        RECT 22.600 176.960 22.920 177.020 ;
        RECT 28.580 176.960 28.900 177.220 ;
        RECT 31.340 176.960 31.660 177.220 ;
        RECT 41.000 176.960 41.320 177.220 ;
        RECT 12.905 176.820 13.195 176.865 ;
        RECT 14.795 176.820 15.085 176.865 ;
        RECT 17.915 176.820 18.205 176.865 ;
        RECT 12.905 176.680 18.205 176.820 ;
        RECT 12.905 176.635 13.195 176.680 ;
        RECT 14.795 176.635 15.085 176.680 ;
        RECT 17.915 176.635 18.205 176.680 ;
        RECT 20.775 176.635 21.065 176.865 ;
        RECT 28.670 176.820 28.810 176.960 ;
        RECT 31.430 176.820 31.570 176.960 ;
        RECT 35.940 176.820 36.260 176.880 ;
        RECT 41.090 176.820 41.230 176.960 ;
        RECT 22.690 176.680 28.810 176.820 ;
        RECT 30.810 176.680 31.570 176.820 ;
        RECT 31.890 176.680 41.230 176.820 ;
        RECT 12.035 176.480 12.325 176.525 ;
        RECT 13.860 176.480 14.180 176.540 ;
        RECT 12.035 176.340 14.180 176.480 ;
        RECT 12.035 176.295 12.325 176.340 ;
        RECT 13.860 176.280 14.180 176.340 ;
        RECT 17.080 176.480 17.400 176.540 ;
        RECT 17.080 176.340 19.150 176.480 ;
        RECT 17.080 176.280 17.400 176.340 ;
        RECT 19.010 176.200 19.150 176.340 ;
        RECT 12.500 176.140 12.790 176.185 ;
        RECT 14.335 176.140 14.625 176.185 ;
        RECT 17.915 176.140 18.205 176.185 ;
        RECT 12.500 176.000 18.205 176.140 ;
        RECT 12.500 175.955 12.790 176.000 ;
        RECT 14.335 175.955 14.625 176.000 ;
        RECT 17.915 175.955 18.205 176.000 ;
        RECT 18.920 176.160 19.240 176.200 ;
        RECT 18.920 175.940 19.285 176.160 ;
        RECT 19.840 175.940 20.160 176.200 ;
        RECT 18.995 175.845 19.285 175.940 ;
        RECT 13.415 175.615 13.705 175.845 ;
        RECT 15.695 175.800 16.345 175.845 ;
        RECT 18.995 175.800 19.585 175.845 ;
        RECT 15.695 175.660 19.585 175.800 ;
        RECT 15.695 175.615 16.345 175.660 ;
        RECT 19.295 175.615 19.585 175.660 ;
        RECT 13.490 175.460 13.630 175.615 ;
        RECT 14.320 175.460 14.640 175.520 ;
        RECT 13.490 175.320 14.640 175.460 ;
        RECT 19.930 175.460 20.070 175.940 ;
        RECT 20.850 175.800 20.990 176.635 ;
        RECT 22.690 176.185 22.830 176.680 ;
        RECT 23.535 176.480 23.825 176.525 ;
        RECT 23.980 176.480 24.300 176.540 ;
        RECT 23.535 176.340 24.300 176.480 ;
        RECT 23.535 176.295 23.825 176.340 ;
        RECT 23.980 176.280 24.300 176.340 ;
        RECT 22.615 175.955 22.905 176.185 ;
        RECT 23.060 176.140 23.380 176.200 ;
        RECT 24.455 176.140 24.745 176.185 ;
        RECT 23.060 176.000 24.745 176.140 ;
        RECT 23.060 175.940 23.380 176.000 ;
        RECT 24.455 175.955 24.745 176.000 ;
        RECT 26.740 175.940 27.060 176.200 ;
        RECT 30.810 176.185 30.950 176.680 ;
        RECT 31.355 176.480 31.645 176.525 ;
        RECT 31.890 176.480 32.030 176.680 ;
        RECT 35.940 176.620 36.260 176.680 ;
        RECT 31.355 176.340 32.030 176.480 ;
        RECT 32.350 176.340 35.250 176.480 ;
        RECT 31.355 176.295 31.645 176.340 ;
        RECT 28.595 175.955 28.885 176.185 ;
        RECT 30.735 175.955 31.025 176.185 ;
        RECT 31.800 176.140 32.120 176.200 ;
        RECT 32.350 176.140 32.490 176.340 ;
        RECT 31.800 176.000 32.490 176.140 ;
        RECT 35.110 176.140 35.250 176.340 ;
        RECT 36.860 176.140 37.180 176.200 ;
        RECT 35.110 176.000 37.180 176.140 ;
        RECT 25.820 175.800 26.140 175.860 ;
        RECT 20.850 175.660 26.140 175.800 ;
        RECT 25.820 175.600 26.140 175.660 ;
        RECT 26.295 175.800 26.585 175.845 ;
        RECT 27.660 175.800 27.980 175.860 ;
        RECT 26.295 175.660 27.980 175.800 ;
        RECT 28.670 175.800 28.810 175.955 ;
        RECT 31.800 175.940 32.120 176.000 ;
        RECT 36.860 175.940 37.180 176.000 ;
        RECT 37.320 176.140 37.640 176.200 ;
        RECT 37.795 176.140 38.085 176.185 ;
        RECT 37.320 176.000 38.085 176.140 ;
        RECT 37.320 175.940 37.640 176.000 ;
        RECT 37.795 175.955 38.085 176.000 ;
        RECT 34.560 175.800 34.880 175.860 ;
        RECT 28.670 175.660 34.880 175.800 ;
        RECT 26.295 175.615 26.585 175.660 ;
        RECT 27.660 175.600 27.980 175.660 ;
        RECT 34.560 175.600 34.880 175.660 ;
        RECT 35.035 175.615 35.325 175.845 ;
        RECT 29.515 175.460 29.805 175.505 ;
        RECT 19.930 175.320 29.805 175.460 ;
        RECT 14.320 175.260 14.640 175.320 ;
        RECT 29.515 175.275 29.805 175.320 ;
        RECT 29.960 175.460 30.280 175.520 ;
        RECT 35.110 175.460 35.250 175.615 ;
        RECT 29.960 175.320 35.250 175.460 ;
        RECT 36.860 175.460 37.180 175.520 ;
        RECT 38.255 175.460 38.545 175.505 ;
        RECT 36.860 175.320 38.545 175.460 ;
        RECT 29.960 175.260 30.280 175.320 ;
        RECT 36.860 175.260 37.180 175.320 ;
        RECT 38.255 175.275 38.545 175.320 ;
        RECT 8.270 174.640 43.230 175.120 ;
        RECT 52.350 174.650 52.650 174.680 ;
        RECT 47.820 174.350 52.650 174.650 ;
        RECT 52.350 174.320 52.650 174.350 ;
        RECT 18.920 174.100 19.240 174.160 ;
        RECT 26.740 174.100 27.060 174.160 ;
        RECT 18.920 173.960 27.060 174.100 ;
        RECT 18.920 173.900 19.240 173.960 ;
        RECT 26.740 173.900 27.060 173.960 ;
        RECT 47.775 168.530 48.125 168.560 ;
        RECT 55.245 168.530 55.595 187.860 ;
        RECT 58.510 187.805 59.890 187.860 ;
        RECT 60.700 187.830 60.930 189.720 ;
        RECT 60.440 187.720 60.930 187.830 ;
        RECT 61.340 187.830 61.570 189.720 ;
        RECT 61.340 187.720 61.700 187.830 ;
        RECT 60.440 187.670 60.900 187.720 ;
        RECT 61.370 187.670 61.700 187.720 ;
        RECT 60.440 187.495 60.600 187.670 ;
        RECT 60.390 187.175 60.650 187.495 ;
        RECT 60.980 187.285 61.290 187.515 ;
        RECT 59.775 186.870 60.005 186.930 ;
        RECT 61.085 186.870 61.255 187.285 ;
        RECT 59.775 186.700 61.255 186.870 ;
        RECT 57.570 186.645 58.445 186.665 ;
        RECT 57.570 186.365 58.580 186.645 ;
        RECT 59.775 186.640 60.005 186.700 ;
        RECT 58.340 186.345 58.580 186.365 ;
        RECT 61.540 186.610 61.700 187.670 ;
        RECT 62.105 186.610 62.365 186.690 ;
        RECT 61.540 186.450 62.365 186.610 ;
        RECT 58.370 185.925 58.550 186.345 ;
        RECT 58.370 185.895 61.270 185.925 ;
        RECT 58.370 185.745 61.290 185.895 ;
        RECT 61.000 185.665 61.290 185.745 ;
        RECT 56.865 185.505 57.175 185.535 ;
        RECT 58.510 185.505 59.890 185.565 ;
        RECT 61.540 185.515 61.700 186.450 ;
        RECT 62.105 186.370 62.365 186.450 ;
        RECT 61.280 185.505 61.700 185.515 ;
        RECT 56.865 185.195 59.890 185.505 ;
        RECT 60.810 185.335 61.040 185.505 ;
        RECT 56.865 185.165 57.175 185.195 ;
        RECT 58.510 185.085 59.890 185.195 ;
        RECT 60.440 185.175 61.040 185.335 ;
        RECT 60.440 184.885 60.600 185.175 ;
        RECT 60.810 185.085 61.040 185.175 ;
        RECT 61.250 185.355 61.700 185.505 ;
        RECT 61.250 185.085 61.480 185.355 ;
        RECT 60.360 184.625 60.680 184.885 ;
        RECT 60.950 184.595 61.330 184.945 ;
        RECT 47.775 168.180 55.595 168.530 ;
        RECT 47.775 168.150 48.125 168.180 ;
        RECT 50.450 166.950 50.750 166.980 ;
        RECT 43.820 166.650 50.750 166.950 ;
        RECT 50.450 166.620 50.750 166.650 ;
        RECT 56.000 163.450 56.400 163.500 ;
        RECT 47.720 163.150 56.400 163.450 ;
        RECT 56.000 163.100 56.400 163.150 ;
        RECT 56.885 162.535 57.185 162.565 ;
        RECT 56.005 162.235 57.185 162.535 ;
        RECT 56.005 157.145 56.305 162.235 ;
        RECT 56.885 162.205 57.185 162.235 ;
        RECT 59.755 160.425 60.135 160.775 ;
        RECT 57.215 159.590 57.535 159.850 ;
        RECT 57.255 158.815 57.495 159.590 ;
        RECT 57.255 158.480 58.685 158.815 ;
        RECT 57.305 158.335 58.685 158.480 ;
        RECT 59.495 158.360 59.725 160.250 ;
        RECT 59.235 158.250 59.725 158.360 ;
        RECT 60.135 158.360 60.365 160.250 ;
        RECT 60.135 158.250 60.495 158.360 ;
        RECT 59.235 158.200 59.695 158.250 ;
        RECT 60.165 158.200 60.495 158.250 ;
        RECT 59.235 158.025 59.395 158.200 ;
        RECT 59.185 157.705 59.445 158.025 ;
        RECT 59.775 157.815 60.085 158.045 ;
        RECT 58.570 157.400 58.800 157.460 ;
        RECT 59.880 157.400 60.050 157.815 ;
        RECT 58.570 157.230 60.050 157.400 ;
        RECT 57.135 157.145 57.375 157.175 ;
        RECT 58.570 157.170 58.800 157.230 ;
        RECT 56.005 156.875 57.375 157.145 ;
        RECT 60.335 157.100 60.495 158.200 ;
        RECT 61.415 157.100 61.675 157.180 ;
        RECT 60.335 156.940 61.675 157.100 ;
        RECT 56.005 156.845 57.345 156.875 ;
        RECT 57.165 156.455 57.345 156.845 ;
        RECT 57.165 156.425 60.065 156.455 ;
        RECT 57.165 156.275 60.085 156.425 ;
        RECT 59.795 156.195 60.085 156.275 ;
        RECT 57.305 156.005 58.685 156.095 ;
        RECT 60.335 156.045 60.495 156.940 ;
        RECT 61.415 156.860 61.675 156.940 ;
        RECT 60.075 156.035 60.495 156.045 ;
        RECT 56.710 155.685 58.685 156.005 ;
        RECT 59.605 155.865 59.835 156.035 ;
        RECT 57.305 155.615 58.685 155.685 ;
        RECT 59.235 155.705 59.835 155.865 ;
        RECT 59.235 155.415 59.395 155.705 ;
        RECT 59.605 155.615 59.835 155.705 ;
        RECT 60.045 155.885 60.495 156.035 ;
        RECT 60.045 155.615 60.275 155.885 ;
        RECT 59.155 155.155 59.475 155.415 ;
        RECT 59.745 155.125 60.125 155.475 ;
        RECT 47.720 133.440 58.185 133.765 ;
        RECT 56.930 132.670 57.230 132.700 ;
        RECT 56.075 132.370 57.230 132.670 ;
        RECT 56.075 127.320 56.375 132.370 ;
        RECT 56.930 132.340 57.230 132.370 ;
        RECT 57.860 130.200 58.185 133.440 ;
        RECT 59.590 130.595 59.970 130.945 ;
        RECT 57.050 129.875 58.185 130.200 ;
        RECT 57.050 128.985 57.375 129.875 ;
        RECT 57.050 128.605 58.520 128.985 ;
        RECT 57.140 128.505 58.520 128.605 ;
        RECT 59.330 128.530 59.560 130.420 ;
        RECT 59.070 128.420 59.560 128.530 ;
        RECT 59.970 128.530 60.200 130.420 ;
        RECT 59.970 128.420 60.330 128.530 ;
        RECT 59.070 128.370 59.530 128.420 ;
        RECT 60.000 128.370 60.330 128.420 ;
        RECT 59.070 128.195 59.230 128.370 ;
        RECT 59.020 127.875 59.280 128.195 ;
        RECT 59.610 127.985 59.920 128.215 ;
        RECT 58.405 127.570 58.635 127.630 ;
        RECT 59.715 127.570 59.885 127.985 ;
        RECT 58.405 127.400 59.885 127.570 ;
        RECT 56.970 127.320 57.210 127.345 ;
        RECT 58.405 127.340 58.635 127.400 ;
        RECT 56.075 127.045 57.210 127.320 ;
        RECT 60.170 127.165 60.330 128.370 ;
        RECT 61.290 127.165 61.550 127.245 ;
        RECT 56.075 127.020 57.180 127.045 ;
        RECT 57.000 126.625 57.180 127.020 ;
        RECT 60.170 127.005 61.550 127.165 ;
        RECT 57.000 126.595 59.900 126.625 ;
        RECT 57.000 126.445 59.920 126.595 ;
        RECT 59.630 126.365 59.920 126.445 ;
        RECT 47.780 126.160 48.070 126.190 ;
        RECT 57.140 126.160 58.520 126.265 ;
        RECT 60.170 126.215 60.330 127.005 ;
        RECT 61.290 126.925 61.550 127.005 ;
        RECT 59.910 126.205 60.330 126.215 ;
        RECT 47.780 125.870 58.520 126.160 ;
        RECT 59.440 126.035 59.670 126.205 ;
        RECT 47.780 125.840 48.070 125.870 ;
        RECT 57.140 125.785 58.520 125.870 ;
        RECT 59.070 125.875 59.670 126.035 ;
        RECT 59.070 125.585 59.230 125.875 ;
        RECT 59.440 125.785 59.670 125.875 ;
        RECT 59.880 126.055 60.330 126.205 ;
        RECT 59.880 125.785 60.110 126.055 ;
        RECT 58.990 125.325 59.310 125.585 ;
        RECT 59.580 125.295 59.960 125.645 ;
        RECT 35.825 113.980 36.350 114.445 ;
        RECT 35.855 113.620 36.320 113.980 ;
        RECT 35.850 113.360 36.320 113.620 ;
        RECT 40.800 113.390 41.265 114.485 ;
        RECT 20.700 103.990 21.080 104.340 ;
        RECT 18.250 102.340 19.630 102.380 ;
        RECT 9.980 101.955 19.630 102.340 ;
        RECT 18.250 101.900 19.630 101.955 ;
        RECT 20.440 101.925 20.670 103.815 ;
        RECT 20.180 101.815 20.670 101.925 ;
        RECT 21.080 101.925 21.310 103.815 ;
        RECT 35.850 102.530 36.230 113.360 ;
        RECT 35.390 102.025 35.690 102.385 ;
        RECT 35.830 102.300 36.250 102.530 ;
        RECT 40.865 102.520 41.190 113.390 ;
        RECT 45.765 104.550 46.290 105.015 ;
        RECT 40.865 102.440 41.290 102.520 ;
        RECT 21.080 101.815 21.440 101.925 ;
        RECT 35.830 101.860 36.250 102.090 ;
        RECT 36.400 102.070 37.855 102.370 ;
        RECT 36.410 102.050 36.640 102.070 ;
        RECT 40.425 102.010 40.725 102.370 ;
        RECT 40.870 102.290 41.290 102.440 ;
        RECT 45.795 102.415 46.260 104.550 ;
        RECT 43.405 102.375 43.705 102.405 ;
        RECT 41.460 102.330 43.705 102.375 ;
        RECT 20.180 101.765 20.640 101.815 ;
        RECT 21.110 101.765 21.440 101.815 ;
        RECT 20.180 101.590 20.340 101.765 ;
        RECT 20.130 101.270 20.390 101.590 ;
        RECT 20.720 101.380 21.030 101.610 ;
        RECT 19.515 100.965 19.745 101.025 ;
        RECT 20.825 100.965 20.995 101.380 ;
        RECT 19.515 100.795 20.995 100.965 ;
        RECT 18.080 100.440 18.320 100.740 ;
        RECT 19.515 100.735 19.745 100.795 ;
        RECT 21.280 100.665 21.440 101.765 ;
        RECT 32.790 101.525 33.110 101.535 ;
        RECT 33.805 101.525 34.105 101.585 ;
        RECT 32.790 101.285 34.105 101.525 ;
        RECT 32.790 101.275 33.110 101.285 ;
        RECT 33.805 101.225 34.105 101.285 ;
        RECT 21.250 100.440 24.145 100.665 ;
        RECT 35.875 100.540 36.220 101.860 ;
        RECT 40.870 101.850 41.290 102.080 ;
        RECT 41.450 102.075 43.705 102.330 ;
        RECT 41.450 102.040 41.680 102.075 ;
        RECT 43.405 102.045 43.705 102.075 ;
        RECT 45.375 101.980 45.675 102.340 ;
        RECT 45.830 102.280 46.250 102.415 ;
        RECT 48.090 102.335 48.390 102.365 ;
        RECT 38.525 100.925 38.815 101.155 ;
        RECT 38.585 100.670 38.755 100.925 ;
        RECT 17.275 100.135 17.575 100.165 ;
        RECT 18.110 100.135 18.290 100.440 ;
        RECT 17.275 100.020 18.290 100.135 ;
        RECT 17.275 99.990 21.010 100.020 ;
        RECT 17.275 99.840 21.030 99.990 ;
        RECT 17.275 99.835 18.270 99.840 ;
        RECT 17.275 99.805 17.575 99.835 ;
        RECT 20.740 99.760 21.030 99.840 ;
        RECT 18.250 99.180 19.630 99.660 ;
        RECT 21.280 99.610 21.440 100.440 ;
        RECT 21.020 99.600 21.440 99.610 ;
        RECT 20.550 99.430 20.780 99.600 ;
        RECT 20.180 99.270 20.780 99.430 ;
        RECT 20.180 98.980 20.340 99.270 ;
        RECT 20.550 99.180 20.780 99.270 ;
        RECT 20.990 99.450 21.440 99.600 ;
        RECT 20.990 99.180 21.220 99.450 ;
        RECT 20.100 98.720 20.420 98.980 ;
        RECT 20.690 98.690 21.070 99.040 ;
        RECT 21.530 97.640 21.820 97.870 ;
        RECT 21.590 97.220 21.760 97.640 ;
        RECT 21.545 96.900 21.805 97.220 ;
        RECT 23.920 93.735 24.145 100.440 ;
        RECT 38.540 100.350 38.800 100.670 ;
        RECT 40.890 100.570 41.235 101.850 ;
        RECT 45.830 101.840 46.250 102.070 ;
        RECT 46.400 102.035 48.390 102.335 ;
        RECT 46.410 102.030 46.640 102.035 ;
        RECT 48.090 102.005 48.390 102.035 ;
        RECT 43.280 100.890 43.570 101.120 ;
        RECT 43.340 100.625 43.510 100.890 ;
        RECT 43.295 100.305 43.555 100.625 ;
        RECT 45.880 100.555 46.225 101.840 ;
        RECT 60.050 99.735 60.430 100.085 ;
        RECT 57.600 98.020 58.980 98.125 ;
        RECT 54.740 97.720 58.980 98.020 ;
        RECT 57.600 97.645 58.980 97.720 ;
        RECT 59.790 97.670 60.020 99.560 ;
        RECT 59.530 97.560 60.020 97.670 ;
        RECT 60.430 97.670 60.660 99.560 ;
        RECT 60.430 97.560 60.790 97.670 ;
        RECT 59.530 97.510 59.990 97.560 ;
        RECT 60.460 97.510 60.790 97.560 ;
        RECT 59.530 97.335 59.690 97.510 ;
        RECT 59.480 97.015 59.740 97.335 ;
        RECT 60.070 97.125 60.380 97.355 ;
        RECT 58.865 96.710 59.095 96.770 ;
        RECT 60.175 96.710 60.345 97.125 ;
        RECT 58.865 96.540 60.345 96.710 ;
        RECT 56.005 96.485 57.525 96.505 ;
        RECT 56.005 96.205 57.670 96.485 ;
        RECT 58.865 96.480 59.095 96.540 ;
        RECT 57.430 96.185 57.670 96.205 ;
        RECT 60.630 96.470 60.790 97.510 ;
        RECT 61.755 96.470 62.015 96.550 ;
        RECT 60.630 96.310 62.015 96.470 ;
        RECT 57.460 95.765 57.640 96.185 ;
        RECT 57.460 95.735 60.360 95.765 ;
        RECT 57.460 95.585 60.380 95.735 ;
        RECT 60.090 95.505 60.380 95.585 ;
        RECT 57.600 95.300 58.980 95.405 ;
        RECT 60.630 95.355 60.790 96.310 ;
        RECT 61.755 96.230 62.015 96.310 ;
        RECT 60.370 95.345 60.790 95.355 ;
        RECT 55.895 95.005 58.980 95.300 ;
        RECT 59.900 95.175 60.130 95.345 ;
        RECT 57.600 94.925 58.980 95.005 ;
        RECT 59.530 95.015 60.130 95.175 ;
        RECT 59.530 94.725 59.690 95.015 ;
        RECT 59.900 94.925 60.130 95.015 ;
        RECT 60.340 95.195 60.790 95.345 ;
        RECT 60.340 94.925 60.570 95.195 ;
        RECT 59.450 94.465 59.770 94.725 ;
        RECT 60.040 94.435 60.420 94.785 ;
        RECT 26.020 93.735 26.340 93.755 ;
        RECT 23.920 93.510 26.340 93.735 ;
        RECT 26.020 93.495 26.340 93.510 ;
        RECT 20.850 92.920 21.230 93.270 ;
        RECT 18.400 91.220 19.780 91.310 ;
        RECT 10.125 90.920 19.780 91.220 ;
        RECT 18.400 90.830 19.780 90.920 ;
        RECT 20.590 90.855 20.820 92.745 ;
        RECT 20.330 90.745 20.820 90.855 ;
        RECT 21.230 90.855 21.460 92.745 ;
        RECT 21.230 90.745 21.590 90.855 ;
        RECT 20.330 90.695 20.790 90.745 ;
        RECT 21.260 90.695 21.590 90.745 ;
        RECT 20.330 90.520 20.490 90.695 ;
        RECT 20.280 90.200 20.540 90.520 ;
        RECT 20.870 90.310 21.180 90.540 ;
        RECT 19.665 89.895 19.895 89.955 ;
        RECT 20.975 89.895 21.145 90.310 ;
        RECT 19.665 89.725 21.145 89.895 ;
        RECT 18.230 89.370 18.470 89.670 ;
        RECT 19.665 89.665 19.895 89.725 ;
        RECT 21.430 89.540 21.590 90.695 ;
        RECT 25.895 89.540 26.215 89.560 ;
        RECT 16.145 89.035 16.445 89.065 ;
        RECT 18.260 89.035 18.440 89.370 ;
        RECT 21.400 89.320 26.215 89.540 ;
        RECT 16.145 88.950 18.440 89.035 ;
        RECT 16.145 88.920 21.160 88.950 ;
        RECT 16.145 88.770 21.180 88.920 ;
        RECT 16.145 88.735 18.405 88.770 ;
        RECT 16.145 88.705 16.445 88.735 ;
        RECT 20.890 88.690 21.180 88.770 ;
        RECT 18.400 88.110 19.780 88.590 ;
        RECT 21.430 88.540 21.590 89.320 ;
        RECT 25.895 89.300 26.215 89.320 ;
        RECT 21.170 88.530 21.590 88.540 ;
        RECT 20.700 88.360 20.930 88.530 ;
        RECT 20.330 88.200 20.930 88.360 ;
        RECT 20.330 87.910 20.490 88.200 ;
        RECT 20.700 88.110 20.930 88.200 ;
        RECT 21.140 88.380 21.590 88.530 ;
        RECT 21.140 88.110 21.370 88.380 ;
        RECT 20.250 87.650 20.570 87.910 ;
        RECT 20.840 87.620 21.220 87.970 ;
        RECT 21.665 86.485 21.955 86.715 ;
        RECT 21.725 86.095 21.895 86.485 ;
        RECT 21.680 85.775 21.940 86.095 ;
        RECT 25.985 84.925 26.305 84.950 ;
        RECT 24.115 84.710 26.305 84.925 ;
        RECT 20.800 81.790 21.180 82.140 ;
        RECT 18.350 80.065 19.730 80.180 ;
        RECT 9.835 79.795 19.730 80.065 ;
        RECT 18.350 79.700 19.730 79.795 ;
        RECT 20.540 79.725 20.770 81.615 ;
        RECT 20.280 79.615 20.770 79.725 ;
        RECT 21.180 79.725 21.410 81.615 ;
        RECT 21.180 79.615 21.540 79.725 ;
        RECT 20.280 79.565 20.740 79.615 ;
        RECT 21.210 79.565 21.540 79.615 ;
        RECT 20.280 79.390 20.440 79.565 ;
        RECT 20.230 79.070 20.490 79.390 ;
        RECT 20.820 79.180 21.130 79.410 ;
        RECT 19.615 78.765 19.845 78.825 ;
        RECT 20.925 78.765 21.095 79.180 ;
        RECT 19.615 78.595 21.095 78.765 ;
        RECT 18.180 78.240 18.420 78.540 ;
        RECT 19.615 78.535 19.845 78.595 ;
        RECT 21.380 78.505 21.540 79.565 ;
        RECT 24.115 78.505 24.330 84.710 ;
        RECT 25.985 84.690 26.305 84.710 ;
        RECT 34.710 81.375 34.970 81.695 ;
        RECT 40.255 81.475 40.575 81.735 ;
        RECT 30.065 80.315 34.120 80.610 ;
        RECT 27.040 79.000 28.420 79.480 ;
        RECT 30.065 79.190 30.360 80.315 ;
        RECT 34.755 80.085 34.925 81.375 ;
        RECT 34.695 79.855 34.985 80.085 ;
        RECT 29.245 78.710 29.475 79.000 ;
        RECT 29.680 78.960 30.680 79.190 ;
        RECT 30.890 79.000 31.170 79.015 ;
        RECT 21.355 78.290 24.330 78.505 ;
        RECT 15.110 77.935 15.410 77.965 ;
        RECT 18.210 77.935 18.390 78.240 ;
        RECT 15.110 77.820 18.390 77.935 ;
        RECT 15.110 77.790 21.110 77.820 ;
        RECT 15.110 77.640 21.130 77.790 ;
        RECT 15.110 77.635 18.345 77.640 ;
        RECT 15.110 77.605 15.410 77.635 ;
        RECT 20.840 77.560 21.130 77.640 ;
        RECT 18.350 76.980 19.730 77.460 ;
        RECT 21.380 77.410 21.540 78.290 ;
        RECT 28.295 78.075 28.545 78.135 ;
        RECT 29.260 78.075 29.450 78.710 ;
        RECT 29.680 78.520 30.680 78.750 ;
        RECT 30.885 78.710 31.170 79.000 ;
        RECT 34.590 78.945 35.970 79.425 ;
        RECT 37.615 79.135 37.910 80.500 ;
        RECT 40.330 79.690 40.500 81.475 ;
        RECT 40.270 79.460 40.560 79.690 ;
        RECT 30.890 78.695 31.170 78.710 ;
        RECT 36.795 78.655 37.025 78.945 ;
        RECT 37.230 78.905 38.230 79.135 ;
        RECT 38.440 78.945 38.720 78.960 ;
        RECT 41.585 78.945 42.965 79.425 ;
        RECT 44.610 79.135 44.905 80.595 ;
        RECT 25.275 77.875 25.575 77.905 ;
        RECT 28.295 77.885 29.450 78.075 ;
        RECT 25.275 77.820 26.780 77.875 ;
        RECT 26.960 77.820 27.205 77.865 ;
        RECT 28.295 77.825 28.545 77.885 ;
        RECT 25.275 77.605 27.205 77.820 ;
        RECT 25.275 77.575 26.780 77.605 ;
        RECT 25.275 77.545 25.575 77.575 ;
        RECT 26.960 77.560 27.205 77.605 ;
        RECT 30.075 77.595 30.370 78.520 ;
        RECT 35.845 78.020 36.095 78.080 ;
        RECT 36.810 78.020 37.000 78.655 ;
        RECT 37.230 78.465 38.230 78.695 ;
        RECT 38.435 78.655 38.720 78.945 ;
        RECT 43.790 78.655 44.020 78.945 ;
        RECT 44.225 78.905 45.225 79.135 ;
        RECT 45.435 78.945 45.715 78.960 ;
        RECT 38.440 78.640 38.720 78.655 ;
        RECT 35.845 77.830 37.000 78.020 ;
        RECT 33.035 77.790 33.335 77.820 ;
        RECT 33.035 77.765 34.270 77.790 ;
        RECT 34.510 77.765 34.755 77.810 ;
        RECT 35.845 77.770 36.095 77.830 ;
        RECT 21.120 77.400 21.540 77.410 ;
        RECT 20.650 77.230 20.880 77.400 ;
        RECT 20.280 77.070 20.880 77.230 ;
        RECT 20.280 76.780 20.440 77.070 ;
        RECT 20.650 76.980 20.880 77.070 ;
        RECT 21.090 77.250 21.540 77.400 ;
        RECT 21.090 76.980 21.320 77.250 ;
        RECT 20.200 76.520 20.520 76.780 ;
        RECT 20.790 76.490 21.170 76.840 ;
        RECT 23.010 76.500 23.270 76.820 ;
        RECT 22.165 76.340 22.395 76.400 ;
        RECT 23.055 76.340 23.225 76.500 ;
        RECT 22.165 76.170 23.225 76.340 ;
        RECT 27.040 76.280 28.420 76.760 ;
        RECT 30.065 76.745 30.530 77.595 ;
        RECT 33.035 77.550 34.755 77.765 ;
        RECT 37.625 77.570 37.920 78.465 ;
        RECT 42.840 78.020 43.090 78.080 ;
        RECT 43.805 78.020 43.995 78.655 ;
        RECT 44.225 78.465 45.225 78.695 ;
        RECT 45.430 78.655 45.715 78.945 ;
        RECT 45.435 78.640 45.715 78.655 ;
        RECT 44.620 78.055 44.915 78.465 ;
        RECT 42.840 77.830 43.995 78.020 ;
        RECT 40.300 77.740 40.600 77.770 ;
        RECT 41.505 77.765 41.750 77.810 ;
        RECT 42.840 77.770 43.090 77.830 ;
        RECT 41.110 77.740 41.750 77.765 ;
        RECT 44.625 77.760 44.915 78.055 ;
        RECT 33.035 77.490 34.270 77.550 ;
        RECT 34.510 77.505 34.755 77.550 ;
        RECT 33.035 77.460 33.335 77.490 ;
        RECT 37.585 76.915 38.050 77.570 ;
        RECT 40.300 77.550 41.750 77.740 ;
        RECT 40.300 77.440 41.260 77.550 ;
        RECT 41.505 77.505 41.750 77.550 ;
        RECT 44.620 77.470 44.915 77.760 ;
        RECT 40.300 77.410 40.600 77.440 ;
        RECT 30.035 76.280 30.560 76.745 ;
        RECT 22.165 76.110 22.395 76.170 ;
        RECT 28.055 75.045 28.365 76.280 ;
        RECT 34.590 76.225 35.970 76.705 ;
        RECT 37.585 76.450 38.590 76.915 ;
        RECT 34.635 75.045 34.945 76.225 ;
        RECT 28.055 74.735 34.945 75.045 ;
        RECT 35.580 68.580 35.890 76.225 ;
        RECT 38.125 69.705 38.590 76.450 ;
        RECT 41.585 76.590 42.965 76.705 ;
        RECT 41.585 76.280 43.720 76.590 ;
        RECT 41.585 76.225 42.965 76.280 ;
        RECT 38.095 69.240 38.620 69.705 ;
        RECT 41.605 68.580 41.915 76.225 ;
        RECT 35.580 68.270 41.915 68.580 ;
        RECT 44.625 67.800 44.915 77.470 ;
        RECT 59.550 69.970 59.930 70.320 ;
        RECT 57.100 68.270 58.480 68.360 ;
        RECT 54.090 67.965 58.480 68.270 ;
        RECT 57.100 67.880 58.480 67.965 ;
        RECT 59.290 67.905 59.520 69.795 ;
        RECT 27.620 67.510 44.915 67.800 ;
        RECT 59.030 67.795 59.520 67.905 ;
        RECT 59.930 67.905 60.160 69.795 ;
        RECT 59.930 67.795 60.290 67.905 ;
        RECT 59.030 67.745 59.490 67.795 ;
        RECT 59.960 67.745 60.290 67.795 ;
        RECT 59.030 67.570 59.190 67.745 ;
        RECT 58.980 67.250 59.240 67.570 ;
        RECT 59.570 67.360 59.880 67.590 ;
        RECT 58.365 66.945 58.595 67.005 ;
        RECT 59.675 66.945 59.845 67.360 ;
        RECT 58.365 66.775 59.845 66.945 ;
        RECT 55.830 66.720 57.010 66.745 ;
        RECT 55.830 66.445 57.170 66.720 ;
        RECT 58.365 66.715 58.595 66.775 ;
        RECT 56.930 66.420 57.170 66.445 ;
        RECT 60.130 66.675 60.290 67.745 ;
        RECT 61.160 66.675 61.480 66.725 ;
        RECT 60.130 66.515 61.480 66.675 ;
        RECT 56.960 66.000 57.140 66.420 ;
        RECT 56.960 65.970 59.860 66.000 ;
        RECT 56.960 65.820 59.880 65.970 ;
        RECT 59.590 65.740 59.880 65.820 ;
        RECT 57.100 65.585 58.480 65.640 ;
        RECT 60.130 65.590 60.290 66.515 ;
        RECT 61.160 66.465 61.480 66.515 ;
        RECT 55.750 65.295 58.480 65.585 ;
        RECT 59.870 65.580 60.290 65.590 ;
        RECT 59.400 65.410 59.630 65.580 ;
        RECT 57.100 65.160 58.480 65.295 ;
        RECT 59.030 65.250 59.630 65.410 ;
        RECT 59.030 64.960 59.190 65.250 ;
        RECT 59.400 65.160 59.630 65.250 ;
        RECT 59.840 65.430 60.290 65.580 ;
        RECT 59.840 65.160 60.070 65.430 ;
        RECT 58.950 64.700 59.270 64.960 ;
        RECT 59.540 64.670 59.920 65.020 ;
        RECT 59.420 40.475 59.800 40.825 ;
        RECT 56.970 38.795 58.350 38.865 ;
        RECT 54.680 38.470 58.350 38.795 ;
        RECT 56.970 38.385 58.350 38.470 ;
        RECT 59.160 38.410 59.390 40.300 ;
        RECT 58.900 38.300 59.390 38.410 ;
        RECT 59.800 38.410 60.030 40.300 ;
        RECT 59.800 38.300 60.160 38.410 ;
        RECT 58.900 38.250 59.360 38.300 ;
        RECT 59.830 38.250 60.160 38.300 ;
        RECT 58.900 38.075 59.060 38.250 ;
        RECT 58.850 37.755 59.110 38.075 ;
        RECT 59.440 37.865 59.750 38.095 ;
        RECT 58.235 37.450 58.465 37.510 ;
        RECT 59.545 37.450 59.715 37.865 ;
        RECT 58.235 37.280 59.715 37.450 ;
        RECT 56.800 37.200 57.040 37.225 ;
        RECT 58.235 37.220 58.465 37.280 ;
        RECT 55.885 36.925 57.040 37.200 ;
        RECT 60.000 36.940 60.160 38.250 ;
        RECT 61.160 36.940 61.480 36.990 ;
        RECT 55.885 36.900 57.010 36.925 ;
        RECT 56.830 36.505 57.010 36.900 ;
        RECT 60.000 36.780 61.480 36.940 ;
        RECT 56.830 36.475 59.730 36.505 ;
        RECT 56.830 36.325 59.750 36.475 ;
        RECT 59.460 36.245 59.750 36.325 ;
        RECT 56.970 36.075 58.350 36.145 ;
        RECT 60.000 36.095 60.160 36.780 ;
        RECT 61.160 36.730 61.480 36.780 ;
        RECT 59.740 36.085 60.160 36.095 ;
        RECT 55.880 35.770 58.350 36.075 ;
        RECT 59.270 35.915 59.500 36.085 ;
        RECT 56.970 35.665 58.350 35.770 ;
        RECT 58.900 35.755 59.500 35.915 ;
        RECT 58.900 35.465 59.060 35.755 ;
        RECT 59.270 35.665 59.500 35.755 ;
        RECT 59.710 35.935 60.160 36.085 ;
        RECT 59.710 35.665 59.940 35.935 ;
        RECT 58.820 35.205 59.140 35.465 ;
        RECT 59.410 35.175 59.790 35.525 ;
        RECT 60.450 8.760 60.830 9.110 ;
        RECT 58.000 7.075 59.380 7.150 ;
        RECT 55.855 6.780 59.380 7.075 ;
        RECT 58.000 6.670 59.380 6.780 ;
        RECT 60.190 6.695 60.420 8.585 ;
        RECT 59.930 6.585 60.420 6.695 ;
        RECT 60.830 6.695 61.060 8.585 ;
        RECT 60.830 6.585 61.190 6.695 ;
        RECT 59.930 6.535 60.390 6.585 ;
        RECT 60.860 6.535 61.190 6.585 ;
        RECT 59.930 6.360 60.090 6.535 ;
        RECT 59.880 6.040 60.140 6.360 ;
        RECT 60.470 6.150 60.780 6.380 ;
        RECT 59.265 5.735 59.495 5.795 ;
        RECT 60.575 5.735 60.745 6.150 ;
        RECT 59.265 5.565 60.745 5.735 ;
        RECT 61.030 5.750 61.190 6.535 ;
        RECT 56.845 5.510 58.005 5.555 ;
        RECT 56.845 5.255 58.070 5.510 ;
        RECT 59.265 5.505 59.495 5.565 ;
        RECT 57.830 5.210 58.070 5.255 ;
        RECT 61.030 5.420 62.340 5.750 ;
        RECT 57.860 4.790 58.040 5.210 ;
        RECT 57.860 4.760 60.760 4.790 ;
        RECT 57.860 4.610 60.780 4.760 ;
        RECT 60.490 4.530 60.780 4.610 ;
        RECT 58.000 4.300 59.380 4.430 ;
        RECT 61.030 4.380 61.190 5.420 ;
        RECT 60.770 4.370 61.190 4.380 ;
        RECT 56.805 4.000 59.380 4.300 ;
        RECT 60.300 4.200 60.530 4.370 ;
        RECT 58.000 3.950 59.380 4.000 ;
        RECT 59.930 4.040 60.530 4.200 ;
        RECT 59.930 3.750 60.090 4.040 ;
        RECT 60.300 3.950 60.530 4.040 ;
        RECT 60.740 4.220 61.190 4.370 ;
        RECT 60.740 3.950 60.970 4.220 ;
        RECT 59.850 3.490 60.170 3.750 ;
        RECT 60.440 3.460 60.820 3.810 ;
      LAYER met2 ;
        RECT 46.750 223.840 47.050 223.850 ;
        RECT 46.715 223.560 47.085 223.840 ;
        RECT 33.160 220.750 33.440 220.785 ;
        RECT 31.850 220.740 33.450 220.750 ;
        RECT 6.060 216.740 6.340 220.740 ;
        RECT 15.720 219.550 16.000 220.740 ;
        RECT 15.720 218.640 16.050 219.550 ;
        RECT 15.715 218.360 16.085 218.640 ;
        RECT 15.720 218.350 16.050 218.360 ;
        RECT 15.720 217.450 16.000 218.350 ;
        RECT 15.720 217.310 16.390 217.450 ;
        RECT 15.720 216.740 16.000 217.310 ;
        RECT 6.130 205.470 6.270 216.740 ;
        RECT 16.250 211.330 16.390 217.310 ;
        RECT 22.160 216.740 22.440 220.740 ;
        RECT 31.820 220.450 33.450 220.740 ;
        RECT 31.820 216.740 32.100 220.450 ;
        RECT 33.160 220.415 33.440 220.450 ;
        RECT 41.470 220.355 41.770 220.745 ;
        RECT 41.480 216.740 41.760 220.355 ;
        RECT 46.750 217.905 47.050 223.560 ;
        RECT 121.750 223.285 122.050 223.295 ;
        RECT 62.870 223.140 63.170 223.150 ;
        RECT 70.230 223.140 70.530 223.150 ;
        RECT 73.910 223.140 74.210 223.150 ;
        RECT 59.190 223.040 59.490 223.050 ;
        RECT 48.760 222.950 49.040 222.985 ;
        RECT 47.920 219.450 48.200 220.740 ;
        RECT 47.920 219.150 48.280 219.450 ;
        RECT 47.920 218.350 48.250 219.150 ;
        RECT 47.920 216.740 48.200 218.350 ;
        RECT 16.640 215.410 16.920 215.525 ;
        RECT 16.640 215.270 17.310 215.410 ;
        RECT 16.640 215.155 16.920 215.270 ;
        RECT 16.250 211.190 16.850 211.330 ;
        RECT 10.200 208.355 10.480 208.725 ;
        RECT 16.710 208.530 16.850 211.190 ;
        RECT 6.070 205.150 6.330 205.470 ;
        RECT 10.270 204.450 10.410 208.355 ;
        RECT 16.650 208.210 16.910 208.530 ;
        RECT 15.165 207.335 16.705 207.705 ;
        RECT 17.170 206.830 17.310 215.270 ;
        RECT 17.570 208.210 17.830 208.530 ;
        RECT 17.630 207.170 17.770 208.210 ;
        RECT 17.570 206.850 17.830 207.170 ;
        RECT 17.110 206.510 17.370 206.830 ;
        RECT 11.130 206.170 11.390 206.490 ;
        RECT 13.890 206.170 14.150 206.490 ;
        RECT 18.030 206.170 18.290 206.490 ;
        RECT 10.210 204.130 10.470 204.450 ;
        RECT 11.190 203.430 11.330 206.170 ;
        RECT 11.865 204.615 13.405 204.985 ;
        RECT 13.950 204.450 14.090 206.170 ;
        RECT 15.270 205.150 15.530 205.470 ;
        RECT 13.890 204.130 14.150 204.450 ;
        RECT 14.810 204.130 15.070 204.450 ;
        RECT 14.870 203.430 15.010 204.130 ;
        RECT 15.330 203.770 15.470 205.150 ;
        RECT 15.270 203.450 15.530 203.770 ;
        RECT 11.130 203.110 11.390 203.430 ;
        RECT 13.890 203.110 14.150 203.430 ;
        RECT 14.810 203.110 15.070 203.430 ;
        RECT 16.190 203.285 16.450 203.430 ;
        RECT 10.210 202.770 10.470 203.090 ;
        RECT 11.590 202.770 11.850 203.090 ;
        RECT 9.750 200.730 10.010 201.050 ;
        RECT 7.440 198.155 7.720 198.525 ;
        RECT 7.450 198.010 7.710 198.155 ;
        RECT 8.820 197.475 9.100 197.845 ;
        RECT 8.890 193.570 9.030 197.475 ;
        RECT 9.810 196.290 9.950 200.730 ;
        RECT 10.270 197.900 10.410 202.770 ;
        RECT 11.650 201.730 11.790 202.770 ;
        RECT 11.590 201.410 11.850 201.730 ;
        RECT 11.130 200.730 11.390 201.050 ;
        RECT 10.670 199.710 10.930 200.030 ;
        RECT 10.730 198.670 10.870 199.710 ;
        RECT 10.670 198.350 10.930 198.670 ;
        RECT 10.270 197.760 10.870 197.900 ;
        RECT 10.210 196.990 10.470 197.310 ;
        RECT 9.750 195.970 10.010 196.290 ;
        RECT 9.290 194.610 9.550 194.930 ;
        RECT 8.830 193.250 9.090 193.570 ;
        RECT 7.450 188.830 7.710 189.150 ;
        RECT 4.705 188.050 5.095 188.350 ;
        RECT 7.510 188.325 7.650 188.830 ;
        RECT 2.850 183.390 3.110 183.710 ;
        RECT 2.910 168.000 3.050 183.390 ;
        RECT 3.805 171.050 4.195 171.350 ;
        RECT 2.840 164.000 3.120 168.000 ;
        RECT 3.850 161.550 4.150 171.050 ;
        RECT 4.750 162.450 5.050 188.050 ;
        RECT 7.440 187.955 7.720 188.325 ;
        RECT 8.890 184.730 9.030 193.250 ;
        RECT 9.350 193.230 9.490 194.610 ;
        RECT 9.290 192.910 9.550 193.230 ;
        RECT 9.290 191.890 9.550 192.210 ;
        RECT 9.350 189.830 9.490 191.890 ;
        RECT 9.290 189.510 9.550 189.830 ;
        RECT 9.350 185.410 9.490 189.510 ;
        RECT 9.750 186.450 10.010 186.770 ;
        RECT 9.290 185.090 9.550 185.410 ;
        RECT 8.830 184.410 9.090 184.730 ;
        RECT 5.605 181.150 5.995 181.450 ;
        RECT 5.650 163.450 5.950 181.150 ;
        RECT 9.810 177.870 9.950 186.450 ;
        RECT 10.270 182.690 10.410 196.990 ;
        RECT 10.730 192.890 10.870 197.760 ;
        RECT 11.190 195.610 11.330 200.730 ;
        RECT 11.865 199.175 13.405 199.545 ;
        RECT 11.590 198.690 11.850 199.010 ;
        RECT 11.130 195.290 11.390 195.610 ;
        RECT 11.650 194.500 11.790 198.690 ;
        RECT 13.950 198.410 14.090 203.110 ;
        RECT 16.180 202.915 16.460 203.285 ;
        RECT 17.110 202.770 17.370 203.090 ;
        RECT 14.350 202.430 14.610 202.750 ;
        RECT 14.410 201.050 14.550 202.430 ;
        RECT 15.165 201.895 16.705 202.265 ;
        RECT 14.810 201.410 15.070 201.730 ;
        RECT 14.350 200.730 14.610 201.050 ;
        RECT 14.410 199.010 14.550 200.730 ;
        RECT 14.350 198.690 14.610 199.010 ;
        RECT 13.950 198.270 14.550 198.410 ;
        RECT 13.890 196.990 14.150 197.310 ;
        RECT 13.950 195.805 14.090 196.990 ;
        RECT 13.880 195.435 14.160 195.805 ;
        RECT 13.890 194.950 14.150 195.270 ;
        RECT 13.950 194.590 14.090 194.950 ;
        RECT 11.190 194.360 11.790 194.500 ;
        RECT 10.670 192.570 10.930 192.890 ;
        RECT 11.190 192.550 11.330 194.360 ;
        RECT 13.890 194.270 14.150 194.590 ;
        RECT 11.865 193.735 13.405 194.105 ;
        RECT 14.410 193.480 14.550 198.270 ;
        RECT 14.870 197.990 15.010 201.410 ;
        RECT 15.270 200.390 15.530 200.710 ;
        RECT 15.330 197.990 15.470 200.390 ;
        RECT 16.180 198.835 16.460 199.205 ;
        RECT 16.250 198.330 16.390 198.835 ;
        RECT 16.190 198.010 16.450 198.330 ;
        RECT 14.810 197.670 15.070 197.990 ;
        RECT 15.270 197.670 15.530 197.990 ;
        RECT 16.250 197.845 16.390 198.010 ;
        RECT 14.870 195.690 15.010 197.670 ;
        RECT 16.180 197.475 16.460 197.845 ;
        RECT 15.165 196.455 16.705 196.825 ;
        RECT 17.170 196.290 17.310 202.770 ;
        RECT 17.570 197.670 17.830 197.990 ;
        RECT 17.630 196.370 17.770 197.670 ;
        RECT 18.090 197.310 18.230 206.170 ;
        RECT 22.230 206.150 22.370 216.740 ;
        RECT 25.850 207.870 26.110 208.190 ;
        RECT 29.070 207.870 29.330 208.190 ;
        RECT 23.900 207.335 25.440 207.705 ;
        RECT 22.630 206.850 22.890 207.170 ;
        RECT 22.170 205.830 22.430 206.150 ;
        RECT 18.490 205.490 18.750 205.810 ;
        RECT 18.550 199.205 18.690 205.490 ;
        RECT 20.600 204.615 22.140 204.985 ;
        RECT 19.410 202.430 19.670 202.750 ;
        RECT 18.950 200.390 19.210 200.710 ;
        RECT 18.480 198.835 18.760 199.205 ;
        RECT 18.490 198.350 18.750 198.670 ;
        RECT 18.030 196.990 18.290 197.310 ;
        RECT 17.110 195.970 17.370 196.290 ;
        RECT 17.630 196.230 18.230 196.370 ;
        RECT 14.870 195.550 15.930 195.690 ;
        RECT 13.030 193.340 14.550 193.480 ;
        RECT 13.030 192.550 13.170 193.340 ;
        RECT 15.790 192.970 15.930 195.550 ;
        RECT 16.650 194.950 16.910 195.270 ;
        RECT 16.710 194.330 16.850 194.950 ;
        RECT 18.090 194.930 18.230 196.230 ;
        RECT 18.030 194.610 18.290 194.930 ;
        RECT 16.710 194.190 17.770 194.330 ;
        RECT 13.950 192.890 15.930 192.970 ;
        RECT 17.110 192.910 17.370 193.230 ;
        RECT 13.950 192.830 15.990 192.890 ;
        RECT 11.130 192.230 11.390 192.550 ;
        RECT 12.970 192.230 13.230 192.550 ;
        RECT 11.130 191.550 11.390 191.870 ;
        RECT 12.970 191.550 13.230 191.870 ;
        RECT 10.670 189.850 10.930 190.170 ;
        RECT 10.730 185.410 10.870 189.850 ;
        RECT 11.190 187.110 11.330 191.550 ;
        RECT 13.030 190.510 13.170 191.550 ;
        RECT 13.950 190.850 14.090 192.830 ;
        RECT 15.730 192.570 15.990 192.830 ;
        RECT 14.810 191.550 15.070 191.870 ;
        RECT 13.890 190.530 14.150 190.850 ;
        RECT 12.970 190.190 13.230 190.510 ;
        RECT 13.490 189.430 14.550 189.570 ;
        RECT 13.490 189.150 13.630 189.430 ;
        RECT 13.430 188.830 13.690 189.150 ;
        RECT 13.890 188.830 14.150 189.150 ;
        RECT 11.865 188.295 13.405 188.665 ;
        RECT 13.950 187.450 14.090 188.830 ;
        RECT 13.890 187.130 14.150 187.450 ;
        RECT 11.130 186.790 11.390 187.110 ;
        RECT 12.510 186.450 12.770 186.770 ;
        RECT 12.970 186.450 13.230 186.770 ;
        RECT 10.670 185.090 10.930 185.410 ;
        RECT 10.670 184.070 10.930 184.390 ;
        RECT 11.130 184.070 11.390 184.390 ;
        RECT 10.210 182.370 10.470 182.690 ;
        RECT 10.730 178.950 10.870 184.070 ;
        RECT 11.190 179.970 11.330 184.070 ;
        RECT 12.570 183.710 12.710 186.450 ;
        RECT 13.030 184.730 13.170 186.450 ;
        RECT 12.970 184.410 13.230 184.730 ;
        RECT 13.890 184.070 14.150 184.390 ;
        RECT 12.510 183.390 12.770 183.710 ;
        RECT 11.865 182.855 13.405 183.225 ;
        RECT 13.950 182.010 14.090 184.070 ;
        RECT 13.890 181.690 14.150 182.010 ;
        RECT 11.130 179.650 11.390 179.970 ;
        RECT 12.970 178.970 13.230 179.290 ;
        RECT 10.670 178.630 10.930 178.950 ;
        RECT 13.030 178.690 13.170 178.970 ;
        RECT 13.950 178.950 14.090 181.690 ;
        RECT 13.420 178.690 13.700 178.805 ;
        RECT 13.030 178.550 13.700 178.690 ;
        RECT 13.890 178.630 14.150 178.950 ;
        RECT 13.420 178.435 13.700 178.550 ;
        RECT 9.350 177.730 9.950 177.870 ;
        RECT 9.350 168.000 9.490 177.730 ;
        RECT 11.865 177.415 13.405 177.785 ;
        RECT 13.950 176.570 14.090 178.630 ;
        RECT 13.890 176.250 14.150 176.570 ;
        RECT 14.410 175.550 14.550 189.430 ;
        RECT 14.870 181.330 15.010 191.550 ;
        RECT 15.165 191.015 16.705 191.385 ;
        RECT 15.270 189.850 15.530 190.170 ;
        RECT 16.650 190.080 16.910 190.170 ;
        RECT 17.170 190.080 17.310 192.910 ;
        RECT 16.650 189.940 17.310 190.080 ;
        RECT 16.650 189.850 16.910 189.940 ;
        RECT 15.330 189.490 15.470 189.850 ;
        RECT 16.710 189.685 16.850 189.850 ;
        RECT 15.270 189.170 15.530 189.490 ;
        RECT 16.640 189.315 16.920 189.685 ;
        RECT 17.110 187.470 17.370 187.790 ;
        RECT 15.165 185.575 16.705 185.945 ;
        RECT 17.170 184.810 17.310 187.470 ;
        RECT 16.710 184.670 17.310 184.810 ;
        RECT 16.710 184.390 16.850 184.670 ;
        RECT 17.630 184.390 17.770 194.190 ;
        RECT 18.090 192.550 18.230 194.610 ;
        RECT 18.550 192.550 18.690 198.350 ;
        RECT 19.010 195.950 19.150 200.390 ;
        RECT 18.950 195.630 19.210 195.950 ;
        RECT 19.470 194.590 19.610 202.430 ;
        RECT 21.250 201.070 21.510 201.390 ;
        RECT 21.310 200.710 21.450 201.070 ;
        RECT 21.250 200.390 21.510 200.710 ;
        RECT 22.690 200.030 22.830 206.850 ;
        RECT 25.910 206.490 26.050 207.870 ;
        RECT 29.130 206.830 29.270 207.870 ;
        RECT 31.890 207.170 32.030 216.740 ;
        RECT 38.260 211.755 38.540 212.125 ;
        RECT 32.635 207.335 34.175 207.705 ;
        RECT 38.330 207.170 38.470 211.755 ;
        RECT 41.550 208.610 41.690 216.740 ;
        RECT 47.150 213.150 47.450 213.180 ;
        RECT 45.605 212.850 47.450 213.150 ;
        RECT 47.150 212.820 47.450 212.850 ;
        RECT 47.150 212.050 47.450 212.080 ;
        RECT 46.405 211.750 47.450 212.050 ;
        RECT 47.150 211.720 47.450 211.750 ;
        RECT 41.090 208.470 41.690 208.610 ;
        RECT 30.450 206.850 30.710 207.170 ;
        RECT 31.830 206.850 32.090 207.170 ;
        RECT 38.270 206.850 38.530 207.170 ;
        RECT 29.070 206.510 29.330 206.830 ;
        RECT 23.550 206.170 23.810 206.490 ;
        RECT 25.850 206.170 26.110 206.490 ;
        RECT 27.690 206.170 27.950 206.490 ;
        RECT 28.150 206.170 28.410 206.490 ;
        RECT 23.610 203.430 23.750 206.170 ;
        RECT 25.910 203.430 26.050 206.170 ;
        RECT 26.770 203.790 27.030 204.110 ;
        RECT 23.550 203.110 23.810 203.430 ;
        RECT 25.850 203.110 26.110 203.430 ;
        RECT 26.310 203.110 26.570 203.430 ;
        RECT 23.610 201.730 23.750 203.110 ;
        RECT 23.900 201.895 25.440 202.265 ;
        RECT 23.550 201.410 23.810 201.730 ;
        RECT 26.370 201.390 26.510 203.110 ;
        RECT 26.310 201.070 26.570 201.390 ;
        RECT 23.090 200.730 23.350 201.050 ;
        RECT 22.630 199.710 22.890 200.030 ;
        RECT 20.600 199.175 22.140 199.545 ;
        RECT 19.870 198.010 20.130 198.330 ;
        RECT 20.330 198.010 20.590 198.330 ;
        RECT 19.410 194.270 19.670 194.590 ;
        RECT 18.030 192.230 18.290 192.550 ;
        RECT 18.490 192.230 18.750 192.550 ;
        RECT 18.090 189.830 18.230 192.230 ;
        RECT 18.950 191.550 19.210 191.870 ;
        RECT 18.030 189.510 18.290 189.830 ;
        RECT 18.490 189.170 18.750 189.490 ;
        RECT 18.030 188.830 18.290 189.150 ;
        RECT 18.090 188.130 18.230 188.830 ;
        RECT 18.030 187.810 18.290 188.130 ;
        RECT 18.550 185.490 18.690 189.170 ;
        RECT 19.010 187.110 19.150 191.550 ;
        RECT 19.410 189.850 19.670 190.170 ;
        RECT 18.950 186.790 19.210 187.110 ;
        RECT 18.950 186.110 19.210 186.430 ;
        RECT 18.090 185.350 18.690 185.490 ;
        RECT 16.650 184.070 16.910 184.390 ;
        RECT 17.570 184.070 17.830 184.390 ;
        RECT 17.110 181.690 17.370 182.010 ;
        RECT 14.810 181.010 15.070 181.330 ;
        RECT 15.165 180.135 16.705 180.505 ;
        RECT 14.810 179.650 15.070 179.970 ;
        RECT 14.870 179.370 15.010 179.650 ;
        RECT 14.870 179.230 16.390 179.370 ;
        RECT 16.250 178.610 16.390 179.230 ;
        RECT 16.190 178.290 16.450 178.610 ;
        RECT 17.170 176.570 17.310 181.690 ;
        RECT 18.090 177.870 18.230 185.350 ;
        RECT 19.010 184.130 19.150 186.110 ;
        RECT 18.550 183.990 19.150 184.130 ;
        RECT 18.550 180.990 18.690 183.990 ;
        RECT 19.470 183.710 19.610 189.850 ;
        RECT 19.930 186.340 20.070 198.010 ;
        RECT 20.390 196.290 20.530 198.010 ;
        RECT 22.690 197.310 22.830 199.710 ;
        RECT 22.630 196.990 22.890 197.310 ;
        RECT 20.330 195.970 20.590 196.290 ;
        RECT 22.630 195.970 22.890 196.290 ;
        RECT 20.600 193.735 22.140 194.105 ;
        RECT 22.690 192.550 22.830 195.970 ;
        RECT 23.150 195.950 23.290 200.730 ;
        RECT 23.900 196.455 25.440 196.825 ;
        RECT 26.370 195.950 26.510 201.070 ;
        RECT 23.090 195.630 23.350 195.950 ;
        RECT 26.310 195.630 26.570 195.950 ;
        RECT 23.090 194.950 23.350 195.270 ;
        RECT 25.850 194.950 26.110 195.270 ;
        RECT 23.150 193.570 23.290 194.950 ;
        RECT 23.090 193.250 23.350 193.570 ;
        RECT 22.630 192.230 22.890 192.550 ;
        RECT 22.690 190.850 22.830 192.230 ;
        RECT 23.550 191.890 23.810 192.210 ;
        RECT 23.610 191.610 23.750 191.890 ;
        RECT 23.150 191.470 23.750 191.610 ;
        RECT 22.630 190.530 22.890 190.850 ;
        RECT 20.600 188.295 22.140 188.665 ;
        RECT 22.690 187.450 22.830 190.530 ;
        RECT 22.630 187.130 22.890 187.450 ;
        RECT 19.930 186.200 20.530 186.340 ;
        RECT 19.870 185.090 20.130 185.410 ;
        RECT 19.410 183.390 19.670 183.710 ;
        RECT 18.490 180.670 18.750 180.990 ;
        RECT 19.930 179.970 20.070 185.090 ;
        RECT 20.390 184.245 20.530 186.200 ;
        RECT 22.170 186.110 22.430 186.430 ;
        RECT 20.320 183.875 20.600 184.245 ;
        RECT 22.230 183.710 22.370 186.110 ;
        RECT 22.170 183.390 22.430 183.710 ;
        RECT 20.600 182.855 22.140 183.225 ;
        RECT 23.150 181.670 23.290 191.470 ;
        RECT 23.900 191.015 25.440 191.385 ;
        RECT 25.910 189.570 26.050 194.950 ;
        RECT 26.370 192.210 26.510 195.630 ;
        RECT 26.310 191.890 26.570 192.210 ;
        RECT 25.450 189.430 26.510 189.570 ;
        RECT 23.550 188.830 23.810 189.150 ;
        RECT 23.610 187.790 23.750 188.830 ;
        RECT 23.550 187.470 23.810 187.790 ;
        RECT 25.450 187.110 25.590 189.430 ;
        RECT 25.850 188.830 26.110 189.150 ;
        RECT 25.390 186.790 25.650 187.110 ;
        RECT 25.910 186.770 26.050 188.830 ;
        RECT 25.850 186.450 26.110 186.770 ;
        RECT 23.550 186.110 23.810 186.430 ;
        RECT 21.710 181.350 21.970 181.670 ;
        RECT 23.090 181.350 23.350 181.670 ;
        RECT 20.790 180.670 21.050 180.990 ;
        RECT 19.870 179.650 20.130 179.970 ;
        RECT 20.850 178.950 20.990 180.670 ;
        RECT 21.770 179.880 21.910 181.350 ;
        RECT 22.630 180.730 22.890 180.990 ;
        RECT 22.630 180.670 23.290 180.730 ;
        RECT 22.690 180.590 23.290 180.670 ;
        RECT 21.770 179.740 22.830 179.880 ;
        RECT 19.870 178.630 20.130 178.950 ;
        RECT 20.790 178.630 21.050 178.950 ;
        RECT 18.090 177.730 18.690 177.870 ;
        RECT 17.110 176.250 17.370 176.570 ;
        RECT 14.350 175.230 14.610 175.550 ;
        RECT 15.165 174.695 16.705 175.065 ;
        RECT 18.550 171.325 18.690 177.730 ;
        RECT 19.930 176.230 20.070 178.630 ;
        RECT 20.600 177.415 22.140 177.785 ;
        RECT 22.690 177.250 22.830 179.740 ;
        RECT 22.630 176.930 22.890 177.250 ;
        RECT 23.150 176.230 23.290 180.590 ;
        RECT 23.610 179.630 23.750 186.110 ;
        RECT 23.900 185.575 25.440 185.945 ;
        RECT 24.010 184.750 24.270 185.070 ;
        RECT 24.070 182.010 24.210 184.750 ;
        RECT 24.010 181.690 24.270 182.010 ;
        RECT 23.900 180.135 25.440 180.505 ;
        RECT 25.910 179.630 26.050 186.450 ;
        RECT 26.370 179.970 26.510 189.430 ;
        RECT 26.310 179.650 26.570 179.970 ;
        RECT 23.550 179.310 23.810 179.630 ;
        RECT 25.850 179.310 26.110 179.630 ;
        RECT 24.010 178.290 24.270 178.610 ;
        RECT 23.550 177.950 23.810 178.270 ;
        RECT 18.950 175.910 19.210 176.230 ;
        RECT 19.870 175.910 20.130 176.230 ;
        RECT 23.090 175.910 23.350 176.230 ;
        RECT 19.010 174.190 19.150 175.910 ;
        RECT 18.950 173.870 19.210 174.190 ;
        RECT 18.480 170.955 18.760 171.325 ;
        RECT 19.010 168.350 19.610 168.490 ;
        RECT 19.010 168.000 19.150 168.350 ;
        RECT 9.280 164.000 9.560 168.000 ;
        RECT 18.940 164.000 19.220 168.000 ;
        RECT 19.470 167.925 19.610 168.350 ;
        RECT 23.610 167.925 23.750 177.950 ;
        RECT 24.070 176.570 24.210 178.290 ;
        RECT 26.370 177.870 26.510 179.650 ;
        RECT 25.910 177.730 26.510 177.870 ;
        RECT 26.830 177.870 26.970 203.790 ;
        RECT 27.750 200.710 27.890 206.170 ;
        RECT 27.690 200.390 27.950 200.710 ;
        RECT 27.230 197.670 27.490 197.990 ;
        RECT 27.290 188.130 27.430 197.670 ;
        RECT 28.210 197.650 28.350 206.170 ;
        RECT 30.510 206.150 30.650 206.850 ;
        RECT 34.590 206.510 34.850 206.830 ;
        RECT 31.370 206.170 31.630 206.490 ;
        RECT 30.450 205.830 30.710 206.150 ;
        RECT 28.610 205.150 28.870 205.470 ;
        RECT 28.670 201.730 28.810 205.150 ;
        RECT 29.335 204.615 30.875 204.985 ;
        RECT 29.060 202.915 29.340 203.285 ;
        RECT 28.610 201.410 28.870 201.730 ;
        RECT 29.130 201.050 29.270 202.915 ;
        RECT 30.450 202.430 30.710 202.750 ;
        RECT 30.510 201.390 30.650 202.430 ;
        RECT 30.450 201.070 30.710 201.390 ;
        RECT 29.070 200.730 29.330 201.050 ;
        RECT 28.610 200.390 28.870 200.710 ;
        RECT 28.150 197.330 28.410 197.650 ;
        RECT 27.690 196.990 27.950 197.310 ;
        RECT 27.750 193.570 27.890 196.990 ;
        RECT 28.670 194.590 28.810 200.390 ;
        RECT 31.430 200.370 31.570 206.170 ;
        RECT 34.130 205.490 34.390 205.810 ;
        RECT 34.190 204.450 34.330 205.490 ;
        RECT 34.130 204.130 34.390 204.450 ;
        RECT 31.830 202.430 32.090 202.750 ;
        RECT 31.890 201.050 32.030 202.430 ;
        RECT 32.635 201.895 34.175 202.265 ;
        RECT 34.650 201.050 34.790 206.510 ;
        RECT 36.890 206.170 37.150 206.490 ;
        RECT 40.570 206.170 40.830 206.490 ;
        RECT 35.510 205.830 35.770 206.150 ;
        RECT 35.050 202.770 35.310 203.090 ;
        RECT 35.110 201.730 35.250 202.770 ;
        RECT 35.570 201.730 35.710 205.830 ;
        RECT 36.950 204.450 37.090 206.170 ;
        RECT 38.070 204.615 39.610 204.985 ;
        RECT 36.890 204.130 37.150 204.450 ;
        RECT 37.350 203.450 37.610 203.770 ;
        RECT 36.430 203.110 36.690 203.430 ;
        RECT 35.050 201.410 35.310 201.730 ;
        RECT 35.510 201.410 35.770 201.730 ;
        RECT 31.830 200.730 32.090 201.050 ;
        RECT 34.590 200.730 34.850 201.050 ;
        RECT 35.510 200.730 35.770 201.050 ;
        RECT 35.970 200.730 36.230 201.050 ;
        RECT 31.370 200.050 31.630 200.370 ;
        RECT 29.335 199.175 30.875 199.545 ;
        RECT 31.890 199.010 32.030 200.730 ;
        RECT 32.290 199.710 32.550 200.030 ;
        RECT 31.830 198.690 32.090 199.010 ;
        RECT 29.530 198.010 29.790 198.330 ;
        RECT 29.590 195.610 29.730 198.010 ;
        RECT 30.910 196.990 31.170 197.310 ;
        RECT 31.830 196.990 32.090 197.310 ;
        RECT 29.530 195.290 29.790 195.610 ;
        RECT 28.610 194.270 28.870 194.590 ;
        RECT 30.970 194.500 31.110 196.990 ;
        RECT 30.970 194.360 31.570 194.500 ;
        RECT 29.335 193.735 30.875 194.105 ;
        RECT 27.690 193.480 27.950 193.570 ;
        RECT 27.690 193.340 28.350 193.480 ;
        RECT 27.690 193.250 27.950 193.340 ;
        RECT 27.230 187.810 27.490 188.130 ;
        RECT 28.210 186.850 28.350 193.340 ;
        RECT 28.610 191.550 28.870 191.870 ;
        RECT 27.750 186.710 28.350 186.850 ;
        RECT 27.750 178.950 27.890 186.710 ;
        RECT 28.670 185.070 28.810 191.550 ;
        RECT 29.335 188.295 30.875 188.665 ;
        RECT 30.910 185.320 31.170 185.410 ;
        RECT 31.430 185.320 31.570 194.360 ;
        RECT 31.890 189.150 32.030 196.990 ;
        RECT 32.350 192.210 32.490 199.710 ;
        RECT 32.635 196.455 34.175 196.825 ;
        RECT 34.650 196.200 34.790 200.730 ;
        RECT 35.050 199.710 35.310 200.030 ;
        RECT 33.730 196.060 34.790 196.200 ;
        RECT 33.730 194.590 33.870 196.060 ;
        RECT 35.110 195.610 35.250 199.710 ;
        RECT 34.590 195.290 34.850 195.610 ;
        RECT 35.050 195.290 35.310 195.610 ;
        RECT 34.650 195.125 34.790 195.290 ;
        RECT 34.580 194.755 34.860 195.125 ;
        RECT 33.670 194.270 33.930 194.590 ;
        RECT 32.290 191.890 32.550 192.210 ;
        RECT 33.730 191.870 33.870 194.270 ;
        RECT 33.670 191.550 33.930 191.870 ;
        RECT 32.635 191.015 34.175 191.385 ;
        RECT 34.650 190.850 34.790 194.755 ;
        RECT 35.110 193.570 35.250 195.290 ;
        RECT 35.050 193.250 35.310 193.570 ;
        RECT 34.590 190.530 34.850 190.850 ;
        RECT 32.290 189.170 32.550 189.490 ;
        RECT 31.830 188.830 32.090 189.150 ;
        RECT 31.830 186.110 32.090 186.430 ;
        RECT 30.910 185.180 31.570 185.320 ;
        RECT 30.910 185.090 31.170 185.180 ;
        RECT 28.610 184.750 28.870 185.070 ;
        RECT 28.150 183.390 28.410 183.710 ;
        RECT 27.690 178.630 27.950 178.950 ;
        RECT 26.830 177.730 27.430 177.870 ;
        RECT 24.010 176.250 24.270 176.570 ;
        RECT 25.910 175.890 26.050 177.730 ;
        RECT 26.770 175.910 27.030 176.230 ;
        RECT 27.290 176.085 27.430 177.730 ;
        RECT 25.850 175.570 26.110 175.890 ;
        RECT 23.900 174.695 25.440 175.065 ;
        RECT 26.830 174.190 26.970 175.910 ;
        RECT 27.220 175.715 27.500 176.085 ;
        RECT 27.690 175.570 27.950 175.890 ;
        RECT 26.770 173.870 27.030 174.190 ;
        RECT 27.750 169.850 27.890 175.570 ;
        RECT 28.210 175.460 28.350 183.390 ;
        RECT 28.670 182.010 28.810 184.750 ;
        RECT 29.335 182.855 30.875 183.225 ;
        RECT 28.610 181.690 28.870 182.010 ;
        RECT 31.890 181.330 32.030 186.110 ;
        RECT 32.350 185.410 32.490 189.170 ;
        RECT 34.590 187.130 34.850 187.450 ;
        RECT 32.635 185.575 34.175 185.945 ;
        RECT 34.650 185.410 34.790 187.130 ;
        RECT 32.290 185.090 32.550 185.410 ;
        RECT 34.590 185.090 34.850 185.410 ;
        RECT 35.110 184.390 35.250 193.250 ;
        RECT 35.050 184.070 35.310 184.390 ;
        RECT 35.050 183.390 35.310 183.710 ;
        RECT 34.590 182.370 34.850 182.690 ;
        RECT 31.830 181.010 32.090 181.330 ;
        RECT 32.290 181.010 32.550 181.330 ;
        RECT 29.070 180.670 29.330 180.990 ;
        RECT 29.130 179.290 29.270 180.670 ;
        RECT 32.350 179.970 32.490 181.010 ;
        RECT 32.635 180.135 34.175 180.505 ;
        RECT 34.650 179.970 34.790 182.370 ;
        RECT 35.110 181.330 35.250 183.390 ;
        RECT 35.050 181.010 35.310 181.330 ;
        RECT 32.290 179.650 32.550 179.970 ;
        RECT 34.590 179.650 34.850 179.970 ;
        RECT 29.070 178.970 29.330 179.290 ;
        RECT 31.370 178.970 31.630 179.290 ;
        RECT 28.610 178.630 28.870 178.950 ;
        RECT 28.670 177.250 28.810 178.630 ;
        RECT 29.335 177.415 30.875 177.785 ;
        RECT 31.430 177.250 31.570 178.970 ;
        RECT 31.820 178.435 32.100 178.805 ;
        RECT 28.610 176.930 28.870 177.250 ;
        RECT 31.370 176.930 31.630 177.250 ;
        RECT 31.890 176.230 32.030 178.435 ;
        RECT 31.830 175.910 32.090 176.230 ;
        RECT 34.590 175.800 34.850 175.890 ;
        RECT 35.110 175.800 35.250 181.010 ;
        RECT 35.570 179.630 35.710 200.730 ;
        RECT 36.030 198.330 36.170 200.730 ;
        RECT 36.490 198.330 36.630 203.110 ;
        RECT 37.410 201.050 37.550 203.450 ;
        RECT 38.270 202.770 38.530 203.090 ;
        RECT 37.350 200.960 37.610 201.050 ;
        RECT 36.950 200.820 37.610 200.960 ;
        RECT 35.970 198.010 36.230 198.330 ;
        RECT 36.430 198.010 36.690 198.330 ;
        RECT 35.960 196.795 36.240 197.165 ;
        RECT 36.030 194.930 36.170 196.795 ;
        RECT 35.970 194.610 36.230 194.930 ;
        RECT 35.970 192.800 36.230 192.890 ;
        RECT 36.490 192.800 36.630 198.010 ;
        RECT 36.950 195.610 37.090 200.820 ;
        RECT 37.350 200.730 37.610 200.820 ;
        RECT 37.810 200.730 38.070 201.050 ;
        RECT 37.870 199.940 38.010 200.730 ;
        RECT 38.330 200.030 38.470 202.770 ;
        RECT 40.110 200.730 40.370 201.050 ;
        RECT 37.410 199.800 38.010 199.940 ;
        RECT 37.410 198.920 37.550 199.800 ;
        RECT 38.270 199.710 38.530 200.030 ;
        RECT 38.070 199.175 39.610 199.545 ;
        RECT 40.170 198.920 40.310 200.730 ;
        RECT 37.410 198.780 38.010 198.920 ;
        RECT 37.870 197.165 38.010 198.780 ;
        RECT 38.330 198.780 40.310 198.920 ;
        RECT 37.800 196.795 38.080 197.165 ;
        RECT 38.330 195.950 38.470 198.780 ;
        RECT 40.110 198.010 40.370 198.330 ;
        RECT 38.730 197.560 38.990 197.650 ;
        RECT 38.730 197.420 39.390 197.560 ;
        RECT 38.730 197.330 38.990 197.420 ;
        RECT 38.270 195.860 38.530 195.950 ;
        RECT 38.270 195.720 38.930 195.860 ;
        RECT 38.270 195.630 38.530 195.720 ;
        RECT 36.890 195.290 37.150 195.610 ;
        RECT 37.800 195.010 38.080 195.125 ;
        RECT 38.270 195.010 38.530 195.270 ;
        RECT 37.800 194.950 38.530 195.010 ;
        RECT 36.890 194.610 37.150 194.930 ;
        RECT 37.800 194.870 38.470 194.950 ;
        RECT 37.800 194.755 38.080 194.870 ;
        RECT 35.970 192.660 36.630 192.800 ;
        RECT 35.970 192.570 36.230 192.660 ;
        RECT 35.970 191.550 36.230 191.870 ;
        RECT 35.510 179.310 35.770 179.630 ;
        RECT 36.030 176.910 36.170 191.550 ;
        RECT 36.490 188.130 36.630 192.660 ;
        RECT 36.950 191.870 37.090 194.610 ;
        RECT 38.790 194.590 38.930 195.720 ;
        RECT 39.250 195.010 39.390 197.420 ;
        RECT 39.650 195.860 39.910 195.950 ;
        RECT 40.170 195.860 40.310 198.010 ;
        RECT 39.650 195.720 40.310 195.860 ;
        RECT 39.650 195.630 39.910 195.720 ;
        RECT 39.250 194.870 40.310 195.010 ;
        RECT 37.810 194.500 38.070 194.590 ;
        RECT 37.410 194.360 38.070 194.500 ;
        RECT 36.890 191.550 37.150 191.870 ;
        RECT 36.430 187.810 36.690 188.130 ;
        RECT 36.490 182.010 36.630 187.810 ;
        RECT 36.950 187.450 37.090 191.550 ;
        RECT 36.890 187.130 37.150 187.450 ;
        RECT 36.890 184.070 37.150 184.390 ;
        RECT 36.430 181.690 36.690 182.010 ;
        RECT 36.950 179.630 37.090 184.070 ;
        RECT 36.890 179.310 37.150 179.630 ;
        RECT 36.890 177.950 37.150 178.270 ;
        RECT 35.970 176.590 36.230 176.910 ;
        RECT 36.950 176.230 37.090 177.950 ;
        RECT 37.410 176.230 37.550 194.360 ;
        RECT 37.810 194.270 38.070 194.360 ;
        RECT 38.730 194.270 38.990 194.590 ;
        RECT 38.070 193.735 39.610 194.105 ;
        RECT 39.650 192.910 39.910 193.230 ;
        RECT 39.710 190.170 39.850 192.910 ;
        RECT 40.170 190.850 40.310 194.870 ;
        RECT 40.110 190.530 40.370 190.850 ;
        RECT 39.650 190.080 39.910 190.170 ;
        RECT 39.650 189.940 40.310 190.080 ;
        RECT 39.650 189.850 39.910 189.940 ;
        RECT 38.070 188.295 39.610 188.665 ;
        RECT 40.170 188.040 40.310 189.940 ;
        RECT 39.710 187.900 40.310 188.040 ;
        RECT 39.710 185.070 39.850 187.900 ;
        RECT 40.110 187.130 40.370 187.450 ;
        RECT 40.170 185.410 40.310 187.130 ;
        RECT 40.630 185.410 40.770 206.170 ;
        RECT 41.090 190.510 41.230 208.470 ;
        RECT 41.370 207.335 42.910 207.705 ;
        RECT 47.990 207.170 48.130 216.740 ;
        RECT 47.930 206.850 48.190 207.170 ;
        RECT 43.790 203.110 44.050 203.430 ;
        RECT 43.330 202.430 43.590 202.750 ;
        RECT 41.370 201.895 42.910 202.265 ;
        RECT 43.390 201.925 43.530 202.430 ;
        RECT 43.320 201.555 43.600 201.925 ;
        RECT 41.370 196.455 42.910 196.825 ;
        RECT 43.850 195.270 43.990 203.110 ;
        RECT 41.950 194.610 42.210 194.930 ;
        RECT 43.320 194.755 43.600 195.125 ;
        RECT 43.790 194.950 44.050 195.270 ;
        RECT 47.550 195.050 47.850 195.080 ;
        RECT 41.490 194.270 41.750 194.590 ;
        RECT 41.550 193.230 41.690 194.270 ;
        RECT 41.490 192.910 41.750 193.230 ;
        RECT 42.010 192.550 42.150 194.610 ;
        RECT 43.390 193.570 43.530 194.755 ;
        RECT 43.330 193.250 43.590 193.570 ;
        RECT 41.950 192.230 42.210 192.550 ;
        RECT 41.370 191.015 42.910 191.385 ;
        RECT 41.030 190.190 41.290 190.510 ;
        RECT 43.330 189.850 43.590 190.170 ;
        RECT 41.030 188.830 41.290 189.150 ;
        RECT 40.110 185.090 40.370 185.410 ;
        RECT 40.570 185.090 40.830 185.410 ;
        RECT 39.650 184.750 39.910 185.070 ;
        RECT 39.710 183.620 39.850 184.750 ;
        RECT 41.090 183.710 41.230 188.830 ;
        RECT 41.370 185.575 42.910 185.945 ;
        RECT 43.390 184.925 43.530 189.850 ;
        RECT 43.850 185.070 43.990 194.950 ;
        RECT 46.805 194.750 47.850 195.050 ;
        RECT 47.550 194.720 47.850 194.750 ;
        RECT 44.710 186.450 44.970 186.770 ;
        RECT 41.490 184.410 41.750 184.730 ;
        RECT 43.320 184.555 43.600 184.925 ;
        RECT 43.790 184.750 44.050 185.070 ;
        RECT 39.710 183.480 40.770 183.620 ;
        RECT 38.070 182.855 39.610 183.225 ;
        RECT 40.630 182.690 40.770 183.480 ;
        RECT 41.030 183.390 41.290 183.710 ;
        RECT 40.570 182.370 40.830 182.690 ;
        RECT 40.110 181.010 40.370 181.330 ;
        RECT 38.270 180.670 38.530 180.990 ;
        RECT 38.330 179.290 38.470 180.670 ;
        RECT 40.170 179.970 40.310 181.010 ;
        RECT 40.110 179.650 40.370 179.970 ;
        RECT 40.630 179.630 40.770 182.370 ;
        RECT 41.550 181.330 41.690 184.410 ;
        RECT 41.950 184.070 42.210 184.390 ;
        RECT 42.010 181.330 42.150 184.070 ;
        RECT 41.490 181.010 41.750 181.330 ;
        RECT 41.950 181.010 42.210 181.330 ;
        RECT 41.370 180.135 42.910 180.505 ;
        RECT 40.570 179.310 40.830 179.630 ;
        RECT 38.270 178.970 38.530 179.290 ;
        RECT 41.030 178.970 41.290 179.290 ;
        RECT 38.070 177.415 39.610 177.785 ;
        RECT 41.090 177.250 41.230 178.970 ;
        RECT 41.030 176.930 41.290 177.250 ;
        RECT 36.890 175.910 37.150 176.230 ;
        RECT 37.350 175.910 37.610 176.230 ;
        RECT 34.590 175.660 35.250 175.800 ;
        RECT 34.590 175.570 34.850 175.660 ;
        RECT 29.990 175.460 30.250 175.550 ;
        RECT 28.210 175.320 30.250 175.460 ;
        RECT 29.990 175.230 30.250 175.320 ;
        RECT 36.890 175.230 37.150 175.550 ;
        RECT 32.635 174.695 34.175 175.065 ;
        RECT 27.750 169.710 28.810 169.850 ;
        RECT 28.670 168.000 28.810 169.710 ;
        RECT 35.110 168.350 35.710 168.490 ;
        RECT 35.110 168.000 35.250 168.350 ;
        RECT 19.400 167.555 19.680 167.925 ;
        RECT 23.540 167.555 23.820 167.925 ;
        RECT 27.360 165.950 27.640 165.985 ;
        RECT 28.600 165.950 28.880 168.000 ;
        RECT 27.350 165.650 28.880 165.950 ;
        RECT 27.360 165.615 27.640 165.650 ;
        RECT 28.600 164.000 28.880 165.650 ;
        RECT 35.040 166.950 35.320 168.000 ;
        RECT 35.570 167.810 35.710 168.350 ;
        RECT 36.950 167.810 37.090 175.230 ;
        RECT 41.370 174.695 42.910 175.065 ;
        RECT 44.770 168.000 44.910 186.450 ;
        RECT 47.850 174.650 48.150 174.680 ;
        RECT 47.105 174.350 48.150 174.650 ;
        RECT 47.850 174.320 48.150 174.350 ;
        RECT 46.750 169.940 47.050 169.950 ;
        RECT 46.715 169.660 47.085 169.940 ;
        RECT 35.570 167.670 37.090 167.810 ;
        RECT 43.850 166.950 44.150 166.980 ;
        RECT 35.040 166.650 44.150 166.950 ;
        RECT 35.040 164.000 35.320 166.650 ;
        RECT 43.850 166.620 44.150 166.650 ;
        RECT 44.700 165.950 44.980 168.000 ;
        RECT 46.750 165.950 47.050 169.660 ;
        RECT 47.745 168.180 48.155 168.530 ;
        RECT 44.700 165.650 47.050 165.950 ;
        RECT 44.700 164.000 44.980 165.650 ;
        RECT 47.775 164.670 48.125 168.180 ;
        RECT 47.730 164.320 48.170 164.670 ;
        RECT 47.750 163.450 48.050 163.480 ;
        RECT 5.650 163.150 48.050 163.450 ;
        RECT 47.750 163.120 48.050 163.150 ;
        RECT 48.170 162.475 48.450 162.510 ;
        RECT 47.660 162.450 48.460 162.475 ;
        RECT 48.750 162.450 49.050 222.950 ;
        RECT 59.155 222.760 59.525 223.040 ;
        RECT 62.835 222.860 63.205 223.140 ;
        RECT 66.550 223.040 66.850 223.050 ;
        RECT 59.190 222.450 59.490 222.760 ;
        RECT 58.320 222.150 59.490 222.450 ;
        RECT 62.870 221.650 63.170 222.860 ;
        RECT 66.515 222.760 66.885 223.040 ;
        RECT 70.195 222.860 70.565 223.140 ;
        RECT 73.875 222.860 74.245 223.140 ;
        RECT 77.590 223.040 77.890 223.050 ;
        RECT 81.270 223.040 81.570 223.050 ;
        RECT 49.750 221.600 63.170 221.650 ;
        RECT 49.600 221.350 63.170 221.600 ;
        RECT 49.600 162.475 49.900 221.350 ;
        RECT 66.550 220.550 66.850 222.760 ;
        RECT 50.450 220.250 66.850 220.550 ;
        RECT 50.450 166.950 50.750 220.250 ;
        RECT 70.230 219.450 70.530 222.860 ;
        RECT 51.320 219.150 70.530 219.450 ;
        RECT 50.420 166.650 50.780 166.950 ;
        RECT 4.750 162.175 48.460 162.450 ;
        RECT 4.750 162.150 47.975 162.175 ;
        RECT 48.170 162.140 48.450 162.175 ;
        RECT 48.715 162.150 49.060 162.450 ;
        RECT 49.555 162.175 49.945 162.475 ;
        RECT 49.585 162.150 49.900 162.175 ;
        RECT 48.750 161.550 49.050 162.150 ;
        RECT 3.850 161.250 49.050 161.550 ;
        RECT 47.750 133.765 48.075 133.795 ;
        RECT 46.300 133.440 48.075 133.765 ;
        RECT 47.750 133.410 48.075 133.440 ;
        RECT 47.775 126.850 48.075 127.240 ;
        RECT 47.780 126.160 48.070 126.850 ;
        RECT 47.750 125.870 48.100 126.160 ;
        RECT 40.810 121.620 41.275 121.645 ;
        RECT 40.790 121.205 41.295 121.620 ;
        RECT 35.805 119.960 36.270 119.985 ;
        RECT 35.785 119.545 36.290 119.960 ;
        RECT 35.805 116.485 36.270 119.545 ;
        RECT 40.810 116.485 41.275 121.205 ;
        RECT 35.805 116.000 36.320 116.485 ;
        RECT 35.855 113.950 36.320 116.000 ;
        RECT 40.800 115.970 41.275 116.485 ;
        RECT 40.800 114.455 41.265 115.970 ;
        RECT 40.770 113.990 41.295 114.455 ;
        RECT 48.750 113.205 49.050 161.250 ;
        RECT 11.615 112.905 49.050 113.205 ;
        RECT 10.010 102.340 10.395 102.370 ;
        RECT 8.250 101.955 10.395 102.340 ;
        RECT 10.010 101.925 10.395 101.955 ;
        RECT 10.155 91.220 10.455 91.250 ;
        RECT 8.320 90.920 10.455 91.220 ;
        RECT 10.155 90.890 10.455 90.920 ;
        RECT 8.415 80.065 8.805 80.080 ;
        RECT 9.865 80.065 10.135 80.095 ;
        RECT 8.415 79.795 10.135 80.065 ;
        RECT 8.415 79.780 8.805 79.795 ;
        RECT 9.865 79.765 10.135 79.795 ;
        RECT 11.615 71.750 11.915 112.905 ;
        RECT 49.600 111.735 49.900 162.150 ;
        RECT 12.910 111.435 49.900 111.735 ;
        RECT 12.910 73.375 13.210 111.435 ;
        RECT 50.450 110.480 50.750 166.650 ;
        RECT 13.970 110.180 50.750 110.480 ;
        RECT 13.970 74.610 14.270 110.180 ;
        RECT 51.350 108.975 51.650 219.150 ;
        RECT 73.910 218.450 74.210 222.860 ;
        RECT 77.555 222.760 77.925 223.040 ;
        RECT 81.235 222.760 81.605 223.040 ;
        RECT 121.715 223.005 122.085 223.285 ;
        RECT 84.950 222.840 85.250 222.850 ;
        RECT 52.350 218.150 74.210 218.450 ;
        RECT 52.350 174.650 52.650 218.150 ;
        RECT 77.590 217.450 77.890 222.760 ;
        RECT 53.250 217.150 77.890 217.450 ;
        RECT 53.250 195.050 53.550 217.150 ;
        RECT 81.270 216.450 81.570 222.760 ;
        RECT 84.915 222.560 85.285 222.840 ;
        RECT 54.250 216.150 81.570 216.450 ;
        RECT 54.250 212.050 54.550 216.150 ;
        RECT 84.950 215.550 85.250 222.560 ;
        RECT 55.250 215.250 85.250 215.550 ;
        RECT 55.250 213.150 55.550 215.250 ;
        RECT 121.750 214.310 122.050 223.005 ;
        RECT 56.020 213.950 56.380 214.250 ;
        RECT 56.875 214.010 122.050 214.310 ;
        RECT 55.220 212.850 55.580 213.150 ;
        RECT 54.220 211.750 54.580 212.050 ;
        RECT 53.220 194.750 53.580 195.050 ;
        RECT 52.320 174.350 52.680 174.650 ;
        RECT 15.110 108.675 51.650 108.975 ;
        RECT 15.110 77.935 15.410 108.675 ;
        RECT 52.350 107.645 52.650 174.350 ;
        RECT 16.145 107.345 52.650 107.645 ;
        RECT 16.145 89.035 16.445 107.345 ;
        RECT 53.250 106.375 53.550 194.750 ;
        RECT 17.275 106.075 53.550 106.375 ;
        RECT 17.275 100.135 17.575 106.075 ;
        RECT 20.070 105.625 20.535 105.650 ;
        RECT 20.050 105.210 20.555 105.625 ;
        RECT 20.070 101.220 20.535 105.210 ;
        RECT 45.795 105.015 46.260 105.045 ;
        RECT 45.795 104.550 47.125 105.015 ;
        RECT 45.795 104.520 46.260 104.550 ;
        RECT 54.250 104.195 54.550 211.750 ;
        RECT 37.525 103.895 54.550 104.195 ;
        RECT 37.525 102.040 37.825 103.895 ;
        RECT 55.250 103.125 55.550 212.850 ;
        RECT 43.405 102.825 55.550 103.125 ;
        RECT 43.405 102.375 43.705 102.825 ;
        RECT 43.375 102.075 43.735 102.375 ;
        RECT 56.050 102.335 56.350 213.950 ;
        RECT 56.875 212.975 57.175 214.010 ;
        RECT 57.600 191.390 57.900 191.400 ;
        RECT 57.565 191.110 57.935 191.390 ;
        RECT 57.600 186.335 57.900 191.110 ;
        RECT 60.360 187.205 60.680 187.465 ;
        RECT 56.835 185.195 57.205 185.505 ;
        RECT 56.865 183.260 57.175 185.195 ;
        RECT 60.440 184.915 60.600 187.205 ;
        RECT 62.085 187.170 62.385 187.560 ;
        RECT 62.155 186.660 62.315 187.170 ;
        RECT 62.075 186.400 62.395 186.660 ;
        RECT 60.390 184.870 60.650 184.915 ;
        RECT 56.820 182.950 57.220 183.260 ;
        RECT 58.760 162.535 59.040 162.570 ;
        RECT 56.855 162.235 59.050 162.535 ;
        RECT 58.760 162.200 59.040 162.235 ;
        RECT 60.340 161.250 60.745 184.870 ;
        RECT 57.225 160.605 57.525 160.995 ;
        RECT 60.335 160.835 60.745 161.250 ;
        RECT 57.255 159.880 57.495 160.605 ;
        RECT 57.245 159.560 57.505 159.880 ;
        RECT 60.335 159.735 60.740 160.835 ;
        RECT 59.065 159.330 60.740 159.735 ;
        RECT 59.065 157.995 59.470 159.330 ;
        RECT 59.065 157.735 59.475 157.995 ;
        RECT 56.740 155.065 57.060 156.035 ;
        RECT 56.695 154.745 57.105 155.065 ;
        RECT 57.955 132.670 58.235 132.705 ;
        RECT 56.900 132.370 58.245 132.670 ;
        RECT 57.955 132.335 58.235 132.370 ;
        RECT 59.065 128.165 59.470 157.735 ;
        RECT 61.350 157.310 61.740 157.610 ;
        RECT 61.465 157.150 61.625 157.310 ;
        RECT 61.385 156.890 61.705 157.150 ;
        RECT 58.990 127.905 59.470 128.165 ;
        RECT 59.065 125.615 59.470 127.905 ;
        RECT 61.260 127.165 61.580 127.215 ;
        RECT 61.825 127.165 62.215 127.235 ;
        RECT 61.260 127.005 62.215 127.165 ;
        RECT 61.260 126.955 61.580 127.005 ;
        RECT 61.825 126.935 62.215 127.005 ;
        RECT 59.020 125.295 59.470 125.615 ;
        RECT 48.060 102.035 56.350 102.335 ;
        RECT 22.355 101.525 22.730 101.595 ;
        RECT 32.820 101.525 33.080 101.565 ;
        RECT 22.355 101.285 33.080 101.525 ;
        RECT 17.245 99.835 17.605 100.135 ;
        RECT 20.180 99.010 20.340 101.220 ;
        RECT 20.130 98.690 20.390 99.010 ;
        RECT 21.515 97.145 21.835 97.190 ;
        RECT 22.355 97.145 22.730 101.285 ;
        RECT 32.820 101.245 33.080 101.285 ;
        RECT 59.065 101.540 59.470 125.295 ;
        RECT 56.035 101.045 56.335 101.055 ;
        RECT 35.845 100.570 36.250 100.915 ;
        RECT 35.875 99.540 36.220 100.570 ;
        RECT 38.510 100.380 38.830 100.640 ;
        RECT 40.860 100.600 41.265 100.945 ;
        RECT 38.585 99.900 38.755 100.380 ;
        RECT 38.520 99.510 38.820 99.900 ;
        RECT 40.890 99.715 41.235 100.600 ;
        RECT 43.265 100.335 43.585 100.595 ;
        RECT 45.850 100.585 46.255 100.930 ;
        RECT 56.000 100.765 56.370 101.045 ;
        RECT 43.340 99.940 43.510 100.335 ;
        RECT 43.275 99.550 43.575 99.940 ;
        RECT 45.880 99.790 46.225 100.585 ;
        RECT 54.770 98.020 55.070 98.050 ;
        RECT 53.150 97.720 55.070 98.020 ;
        RECT 54.770 97.690 55.070 97.720 ;
        RECT 21.515 96.975 22.730 97.145 ;
        RECT 21.515 96.930 21.835 96.975 ;
        RECT 20.125 95.100 20.540 95.120 ;
        RECT 20.100 90.490 20.565 95.100 ;
        RECT 20.100 90.230 20.570 90.490 ;
        RECT 20.100 90.210 20.565 90.230 ;
        RECT 16.115 88.735 16.475 89.035 ;
        RECT 20.330 87.940 20.490 90.210 ;
        RECT 20.280 87.620 20.540 87.940 ;
        RECT 21.650 86.020 21.970 86.065 ;
        RECT 22.355 86.020 22.730 96.975 ;
        RECT 56.035 96.175 56.335 100.765 ;
        RECT 59.065 100.755 59.495 101.540 ;
        RECT 59.090 99.355 59.495 100.755 ;
        RECT 59.090 98.950 59.765 99.355 ;
        RECT 59.360 97.305 59.765 98.950 ;
        RECT 59.360 97.045 59.770 97.305 ;
        RECT 61.690 97.280 62.080 97.580 ;
        RECT 54.580 95.300 54.970 95.305 ;
        RECT 55.925 95.300 56.220 95.330 ;
        RECT 54.580 95.005 56.220 95.300 ;
        RECT 55.925 94.975 56.220 95.005 ;
        RECT 26.050 93.740 26.310 93.785 ;
        RECT 27.670 93.740 28.060 93.780 ;
        RECT 26.050 93.515 28.060 93.740 ;
        RECT 26.050 93.465 26.310 93.515 ;
        RECT 27.670 93.480 28.060 93.515 ;
        RECT 25.925 89.540 26.185 89.590 ;
        RECT 27.495 89.540 27.885 89.580 ;
        RECT 25.925 89.320 27.885 89.540 ;
        RECT 25.925 89.270 26.185 89.320 ;
        RECT 27.495 89.280 27.885 89.320 ;
        RECT 21.650 85.850 22.730 86.020 ;
        RECT 21.650 85.805 21.970 85.850 ;
        RECT 20.200 79.100 20.520 79.360 ;
        RECT 15.080 77.635 15.440 77.935 ;
        RECT 20.280 76.910 20.440 79.100 ;
        RECT 20.175 75.535 20.640 76.910 ;
        RECT 22.355 76.745 22.730 85.850 ;
        RECT 26.015 84.930 26.275 84.980 ;
        RECT 27.655 84.930 28.045 84.975 ;
        RECT 26.015 84.715 28.045 84.930 ;
        RECT 26.015 84.660 26.275 84.715 ;
        RECT 27.655 84.675 28.045 84.715 ;
        RECT 33.795 81.365 34.095 81.755 ;
        RECT 34.680 81.620 35.000 81.665 ;
        RECT 35.605 81.620 35.995 81.685 ;
        RECT 34.680 81.450 35.995 81.620 ;
        RECT 34.680 81.405 35.000 81.450 ;
        RECT 35.605 81.385 35.995 81.450 ;
        RECT 37.615 81.435 37.915 81.825 ;
        RECT 40.285 81.690 40.545 81.765 ;
        RECT 41.545 81.690 41.845 81.800 ;
        RECT 40.285 81.520 41.845 81.690 ;
        RECT 40.285 81.445 40.545 81.520 ;
        RECT 33.795 80.285 34.090 81.365 ;
        RECT 37.615 80.470 37.910 81.435 ;
        RECT 41.545 81.410 41.845 81.520 ;
        RECT 44.610 81.370 44.910 81.760 ;
        RECT 44.610 80.565 44.905 81.370 ;
        RECT 37.585 80.175 37.940 80.470 ;
        RECT 44.580 80.270 44.935 80.565 ;
        RECT 25.245 77.575 25.605 77.875 ;
        RECT 22.980 76.745 23.300 76.790 ;
        RECT 22.355 76.575 23.300 76.745 ;
        RECT 22.355 76.450 22.730 76.575 ;
        RECT 22.980 76.530 23.300 76.575 ;
        RECT 20.200 75.515 20.615 75.535 ;
        RECT 25.275 74.610 25.575 77.575 ;
        RECT 33.005 77.490 33.365 77.790 ;
        RECT 13.970 74.310 25.575 74.610 ;
        RECT 30.065 74.390 30.530 76.775 ;
        RECT 30.045 73.975 30.550 74.390 ;
        RECT 30.065 73.950 30.530 73.975 ;
        RECT 33.035 73.375 33.335 77.490 ;
        RECT 40.270 77.440 40.630 77.740 ;
        RECT 12.910 73.075 33.335 73.375 ;
        RECT 40.300 71.750 40.600 77.440 ;
        RECT 45.670 76.860 46.070 77.170 ;
        RECT 43.380 76.590 43.690 76.620 ;
        RECT 45.715 76.590 46.025 76.860 ;
        RECT 43.380 76.280 46.025 76.590 ;
        RECT 43.380 76.250 43.690 76.280 ;
        RECT 59.360 71.805 59.765 97.045 ;
        RECT 61.805 96.520 61.965 97.280 ;
        RECT 61.725 96.260 62.045 96.520 ;
        RECT 11.615 71.450 40.600 71.750 ;
        RECT 55.860 71.525 56.160 71.535 ;
        RECT 55.825 71.245 56.195 71.525 ;
        RECT 25.100 67.800 25.490 67.805 ;
        RECT 27.650 67.800 27.940 67.830 ;
        RECT 25.100 67.510 27.940 67.800 ;
        RECT 25.100 67.505 25.490 67.510 ;
        RECT 27.650 67.480 27.940 67.510 ;
        RECT 38.125 41.290 38.590 69.735 ;
        RECT 52.660 68.270 52.965 68.315 ;
        RECT 54.120 68.270 54.425 68.300 ;
        RECT 52.660 67.965 54.425 68.270 ;
        RECT 52.660 67.920 52.965 67.965 ;
        RECT 54.120 67.935 54.425 67.965 ;
        RECT 55.860 66.415 56.160 71.245 ;
        RECT 59.350 71.235 59.765 71.805 ;
        RECT 59.350 69.415 59.755 71.235 ;
        RECT 58.825 69.010 59.755 69.415 ;
        RECT 58.825 67.540 59.230 69.010 ;
        RECT 58.825 67.280 59.270 67.540 ;
        RECT 61.795 67.330 62.185 67.630 ;
        RECT 54.175 65.585 54.565 65.590 ;
        RECT 55.780 65.585 56.070 65.615 ;
        RECT 54.175 65.295 56.070 65.585 ;
        RECT 54.175 65.290 54.565 65.295 ;
        RECT 55.780 65.265 56.070 65.295 ;
        RECT 58.825 64.990 59.230 67.280 ;
        RECT 61.190 66.675 61.450 66.755 ;
        RECT 61.910 66.675 62.070 67.330 ;
        RECT 61.190 66.515 62.070 66.675 ;
        RECT 61.190 66.435 61.450 66.515 ;
        RECT 58.825 64.670 59.240 64.990 ;
        RECT 55.925 41.885 56.205 41.920 ;
        RECT 38.105 40.875 38.610 41.290 ;
        RECT 38.125 40.850 38.590 40.875 ;
        RECT 54.710 38.795 55.035 38.825 ;
        RECT 53.375 38.470 55.035 38.795 ;
        RECT 54.710 38.440 55.035 38.470 ;
        RECT 55.915 36.870 56.215 41.885 ;
        RECT 58.825 38.045 59.230 64.670 ;
        RECT 58.820 37.785 59.230 38.045 ;
        RECT 55.910 36.075 56.215 36.105 ;
        RECT 54.320 35.770 56.215 36.075 ;
        RECT 55.910 35.740 56.215 35.770 ;
        RECT 58.825 13.425 59.230 37.785 ;
        RECT 61.775 37.265 62.165 37.565 ;
        RECT 61.190 36.940 61.450 37.020 ;
        RECT 61.890 36.940 62.050 37.265 ;
        RECT 61.190 36.780 62.050 36.940 ;
        RECT 61.190 36.700 61.450 36.780 ;
        RECT 58.825 13.020 60.180 13.425 ;
        RECT 56.875 7.190 57.175 7.200 ;
        RECT 54.555 7.075 54.945 7.080 ;
        RECT 55.885 7.075 56.180 7.105 ;
        RECT 54.555 6.780 56.180 7.075 ;
        RECT 56.840 6.910 57.210 7.190 ;
        RECT 55.885 6.750 56.180 6.780 ;
        RECT 56.875 5.225 57.175 6.910 ;
        RECT 59.775 5.970 60.180 13.020 ;
        RECT 61.980 6.930 62.310 6.955 ;
        RECT 61.960 6.650 62.330 6.930 ;
        RECT 56.835 4.300 57.135 4.330 ;
        RECT 55.685 4.000 57.135 4.300 ;
        RECT 56.835 3.970 57.135 4.000 ;
        RECT 59.930 3.935 60.090 5.970 ;
        RECT 61.980 5.390 62.310 6.650 ;
        RECT 152.575 4.150 153.425 4.170 ;
        RECT 62.430 3.935 153.450 4.150 ;
        RECT 59.825 3.470 153.450 3.935 ;
        RECT 59.880 3.460 60.140 3.470 ;
        RECT 62.430 3.250 153.450 3.470 ;
        RECT 152.575 3.230 153.425 3.250 ;
      LAYER met3 ;
        RECT 46.735 223.850 47.065 223.865 ;
        RECT 51.820 223.850 52.140 223.890 ;
        RECT 40.780 223.750 41.100 223.790 ;
        RECT 1.950 223.450 41.100 223.750 ;
        RECT 46.735 223.550 52.140 223.850 ;
        RECT 55.470 223.640 55.850 223.960 ;
        RECT 59.150 223.640 59.530 223.960 ;
        RECT 62.830 223.740 63.210 224.060 ;
        RECT 66.510 223.740 66.890 224.060 ;
        RECT 70.190 223.740 70.570 224.060 ;
        RECT 46.735 223.535 47.065 223.550 ;
        RECT 51.820 223.510 52.140 223.550 ;
        RECT 1.950 165.950 2.250 223.450 ;
        RECT 40.780 223.410 41.100 223.450 ;
        RECT 4.940 222.950 5.260 222.990 ;
        RECT 3.050 222.650 5.260 222.950 ;
        RECT 3.050 215.640 3.350 222.650 ;
        RECT 4.940 222.610 5.260 222.650 ;
        RECT 48.735 222.950 49.065 222.965 ;
        RECT 55.510 222.950 55.810 223.640 ;
        RECT 59.190 223.065 59.490 223.640 ;
        RECT 62.870 223.165 63.170 223.740 ;
        RECT 48.735 222.650 55.810 222.950 ;
        RECT 59.175 222.735 59.505 223.065 ;
        RECT 62.855 222.835 63.185 223.165 ;
        RECT 66.550 223.065 66.850 223.740 ;
        RECT 70.230 223.165 70.530 223.740 ;
        RECT 73.870 223.640 74.250 223.960 ;
        RECT 77.550 223.740 77.930 224.060 ;
        RECT 73.910 223.165 74.210 223.640 ;
        RECT 66.535 222.735 66.865 223.065 ;
        RECT 70.215 222.835 70.545 223.165 ;
        RECT 73.895 222.835 74.225 223.165 ;
        RECT 77.590 223.065 77.890 223.740 ;
        RECT 81.230 223.540 81.610 223.860 ;
        RECT 84.910 223.640 85.290 223.960 ;
        RECT 121.710 223.745 122.090 224.065 ;
        RECT 81.270 223.065 81.570 223.540 ;
        RECT 77.575 222.735 77.905 223.065 ;
        RECT 81.255 222.735 81.585 223.065 ;
        RECT 84.950 222.865 85.250 223.640 ;
        RECT 121.750 223.310 122.050 223.745 ;
        RECT 121.735 222.980 122.065 223.310 ;
        RECT 48.735 222.635 49.065 222.650 ;
        RECT 84.935 222.535 85.265 222.865 ;
        RECT 154.855 222.010 155.175 222.050 ;
        RECT 41.470 221.710 155.175 222.010 ;
        RECT 33.135 220.750 33.465 220.765 ;
        RECT 40.340 220.750 40.660 220.790 ;
        RECT 33.135 220.450 40.660 220.750 ;
        RECT 41.470 220.725 41.770 221.710 ;
        RECT 154.855 221.670 155.175 221.710 ;
        RECT 33.135 220.435 33.465 220.450 ;
        RECT 40.340 220.410 40.660 220.450 ;
        RECT 41.445 220.375 41.795 220.725 ;
        RECT 112.005 220.420 112.325 220.460 ;
        RECT 104.495 220.120 112.325 220.420 ;
        RECT 15.735 218.650 16.065 218.665 ;
        RECT 15.735 218.350 18.250 218.650 ;
        RECT 15.735 218.335 16.065 218.350 ;
        RECT 2.750 215.490 6.750 215.640 ;
        RECT 16.615 215.490 16.945 215.505 ;
        RECT 2.750 215.190 16.945 215.490 ;
        RECT 2.750 215.040 6.750 215.190 ;
        RECT 16.615 215.175 16.945 215.190 ;
        RECT 17.950 213.150 18.250 218.350 ;
        RECT 46.725 217.925 47.075 218.275 ;
        RECT 46.750 217.090 47.050 217.925 ;
        RECT 46.740 216.710 47.060 217.090 ;
        RECT 57.820 216.425 58.200 216.435 ;
        RECT 104.495 216.425 104.795 220.120 ;
        RECT 112.005 220.080 112.325 220.120 ;
        RECT 112.065 219.620 112.385 219.660 ;
        RECT 57.820 216.125 104.795 216.425 ;
        RECT 105.355 219.320 112.385 219.620 ;
        RECT 57.820 216.115 58.200 216.125 ;
        RECT 58.660 215.360 59.040 215.370 ;
        RECT 105.355 215.360 105.655 219.320 ;
        RECT 112.065 219.280 112.385 219.320 ;
        RECT 106.390 218.765 106.710 218.805 ;
        RECT 112.025 218.765 112.345 218.805 ;
        RECT 106.390 218.465 112.345 218.765 ;
        RECT 106.390 218.425 106.710 218.465 ;
        RECT 112.025 218.425 112.345 218.465 ;
        RECT 107.190 217.715 107.570 217.725 ;
        RECT 111.960 217.715 112.280 217.755 ;
        RECT 107.190 217.415 112.280 217.715 ;
        RECT 107.190 217.405 107.570 217.415 ;
        RECT 111.960 217.375 112.280 217.415 ;
        RECT 108.075 216.445 108.455 216.455 ;
        RECT 111.935 216.445 112.255 216.485 ;
        RECT 108.075 216.145 112.255 216.445 ;
        RECT 108.075 216.135 108.455 216.145 ;
        RECT 111.935 216.105 112.255 216.145 ;
        RECT 58.660 215.060 105.655 215.360 ;
        RECT 108.980 215.295 109.360 215.305 ;
        RECT 111.965 215.295 112.285 215.335 ;
        RECT 58.660 215.050 59.040 215.060 ;
        RECT 108.980 214.995 112.285 215.295 ;
        RECT 108.980 214.985 109.360 214.995 ;
        RECT 111.965 214.955 112.285 214.995 ;
        RECT 51.915 214.505 52.535 214.565 ;
        RECT 112.020 214.505 112.495 214.530 ;
        RECT 51.915 214.020 112.500 214.505 ;
        RECT 51.915 213.580 52.555 214.020 ;
        RECT 112.020 213.995 112.495 214.020 ;
        RECT 45.625 213.150 45.975 213.175 ;
        RECT 17.950 212.850 45.975 213.150 ;
        RECT 45.625 212.825 45.975 212.850 ;
        RECT 38.235 212.090 38.565 212.105 ;
        RECT 44.770 212.090 48.770 212.240 ;
        RECT 38.235 211.790 48.770 212.090 ;
        RECT 38.235 211.775 38.565 211.790 ;
        RECT 44.770 211.640 48.770 211.790 ;
        RECT 2.750 208.690 6.750 208.840 ;
        RECT 10.175 208.690 10.505 208.705 ;
        RECT 2.750 208.390 10.505 208.690 ;
        RECT 2.750 208.240 6.750 208.390 ;
        RECT 10.175 208.375 10.505 208.390 ;
        RECT 15.145 207.355 16.725 207.685 ;
        RECT 23.880 207.355 25.460 207.685 ;
        RECT 32.615 207.355 34.195 207.685 ;
        RECT 41.350 207.355 42.930 207.685 ;
        RECT 11.845 204.635 13.425 204.965 ;
        RECT 20.580 204.635 22.160 204.965 ;
        RECT 29.315 204.635 30.895 204.965 ;
        RECT 38.050 204.635 39.630 204.965 ;
        RECT 16.155 203.250 16.485 203.265 ;
        RECT 29.035 203.250 29.365 203.265 ;
        RECT 16.155 202.950 29.365 203.250 ;
        RECT 16.155 202.935 16.485 202.950 ;
        RECT 29.035 202.935 29.365 202.950 ;
        RECT 15.145 201.915 16.725 202.245 ;
        RECT 23.880 201.915 25.460 202.245 ;
        RECT 32.615 201.915 34.195 202.245 ;
        RECT 41.350 201.915 42.930 202.245 ;
        RECT 43.295 201.890 43.625 201.905 ;
        RECT 44.770 201.890 48.770 202.040 ;
        RECT 43.295 201.590 48.770 201.890 ;
        RECT 43.295 201.575 43.625 201.590 ;
        RECT 44.770 201.440 48.770 201.590 ;
        RECT 4.910 199.740 5.290 200.060 ;
        RECT 4.950 198.640 5.250 199.740 ;
        RECT 11.845 199.195 13.425 199.525 ;
        RECT 20.580 199.195 22.160 199.525 ;
        RECT 29.315 199.195 30.895 199.525 ;
        RECT 38.050 199.195 39.630 199.525 ;
        RECT 16.155 199.170 16.485 199.185 ;
        RECT 18.455 199.170 18.785 199.185 ;
        RECT 16.155 198.870 18.785 199.170 ;
        RECT 16.155 198.855 16.485 198.870 ;
        RECT 18.455 198.855 18.785 198.870 ;
        RECT 2.750 198.490 6.750 198.640 ;
        RECT 7.415 198.490 7.745 198.505 ;
        RECT 2.750 198.190 7.745 198.490 ;
        RECT 2.750 198.040 6.750 198.190 ;
        RECT 7.415 198.175 7.745 198.190 ;
        RECT 8.795 197.810 9.125 197.825 ;
        RECT 16.155 197.810 16.485 197.825 ;
        RECT 8.795 197.510 16.485 197.810 ;
        RECT 8.795 197.495 9.125 197.510 ;
        RECT 16.155 197.495 16.485 197.510 ;
        RECT 35.935 197.130 36.265 197.145 ;
        RECT 37.775 197.130 38.105 197.145 ;
        RECT 35.935 196.830 38.105 197.130 ;
        RECT 35.935 196.815 36.265 196.830 ;
        RECT 37.775 196.815 38.105 196.830 ;
        RECT 15.145 196.475 16.725 196.805 ;
        RECT 23.880 196.475 25.460 196.805 ;
        RECT 32.615 196.475 34.195 196.805 ;
        RECT 41.350 196.475 42.930 196.805 ;
        RECT 13.855 195.780 14.185 195.785 ;
        RECT 13.855 195.770 14.440 195.780 ;
        RECT 13.855 195.470 14.640 195.770 ;
        RECT 13.855 195.460 14.440 195.470 ;
        RECT 13.855 195.455 14.185 195.460 ;
        RECT 34.555 195.090 34.885 195.105 ;
        RECT 37.775 195.090 38.105 195.105 ;
        RECT 34.555 194.790 38.105 195.090 ;
        RECT 34.555 194.775 34.885 194.790 ;
        RECT 37.775 194.775 38.105 194.790 ;
        RECT 43.295 195.090 43.625 195.105 ;
        RECT 44.770 195.090 48.770 195.240 ;
        RECT 43.295 194.790 48.770 195.090 ;
        RECT 43.295 194.775 43.625 194.790 ;
        RECT 44.770 194.640 48.770 194.790 ;
        RECT 11.845 193.755 13.425 194.085 ;
        RECT 20.580 193.755 22.160 194.085 ;
        RECT 29.315 193.755 30.895 194.085 ;
        RECT 38.050 193.755 39.630 194.085 ;
        RECT 15.145 191.035 16.725 191.365 ;
        RECT 23.880 191.035 25.460 191.365 ;
        RECT 32.615 191.035 34.195 191.365 ;
        RECT 41.350 191.035 42.930 191.365 ;
        RECT 16.615 189.650 16.945 189.665 ;
        RECT 17.740 189.650 18.120 189.660 ;
        RECT 16.615 189.350 18.120 189.650 ;
        RECT 16.615 189.335 16.945 189.350 ;
        RECT 17.740 189.340 18.120 189.350 ;
        RECT 2.750 188.290 6.750 188.440 ;
        RECT 11.845 188.315 13.425 188.645 ;
        RECT 20.580 188.315 22.160 188.645 ;
        RECT 29.315 188.315 30.895 188.645 ;
        RECT 38.050 188.315 39.630 188.645 ;
        RECT 7.415 188.290 7.745 188.305 ;
        RECT 2.750 187.990 7.745 188.290 ;
        RECT 2.750 187.840 6.750 187.990 ;
        RECT 7.415 187.975 7.745 187.990 ;
        RECT 15.145 185.595 16.725 185.925 ;
        RECT 23.880 185.595 25.460 185.925 ;
        RECT 32.615 185.595 34.195 185.925 ;
        RECT 41.350 185.595 42.930 185.925 ;
        RECT 51.915 185.040 52.535 213.580 ;
        RECT 56.850 212.995 57.200 213.345 ;
        RECT 56.875 212.240 57.175 212.995 ;
        RECT 56.865 211.860 57.185 212.240 ;
        RECT 63.000 197.230 94.860 213.400 ;
        RECT 43.295 184.890 43.625 184.905 ;
        RECT 44.770 184.890 52.535 185.040 ;
        RECT 43.295 184.590 52.535 184.890 ;
        RECT 43.295 184.575 43.625 184.590 ;
        RECT 44.770 184.440 52.535 184.590 ;
        RECT 51.915 184.430 52.535 184.440 ;
        RECT 53.705 196.765 94.860 197.230 ;
        RECT 20.295 184.210 20.625 184.225 ;
        RECT 16.400 183.910 20.625 184.210 ;
        RECT 11.845 182.875 13.425 183.205 ;
        RECT 2.750 181.490 6.750 181.640 ;
        RECT 16.400 181.490 16.700 183.910 ;
        RECT 20.295 183.895 20.625 183.910 ;
        RECT 20.580 182.875 22.160 183.205 ;
        RECT 29.315 182.875 30.895 183.205 ;
        RECT 38.050 182.875 39.630 183.205 ;
        RECT 2.750 181.190 16.700 181.490 ;
        RECT 2.750 181.040 6.750 181.190 ;
        RECT 15.145 180.155 16.725 180.485 ;
        RECT 23.880 180.155 25.460 180.485 ;
        RECT 32.615 180.155 34.195 180.485 ;
        RECT 41.350 180.155 42.930 180.485 ;
        RECT 13.395 178.770 13.725 178.785 ;
        RECT 17.740 178.770 18.120 178.780 ;
        RECT 31.795 178.770 32.125 178.785 ;
        RECT 13.395 178.470 32.125 178.770 ;
        RECT 13.395 178.455 13.725 178.470 ;
        RECT 17.740 178.460 18.120 178.470 ;
        RECT 31.795 178.455 32.125 178.470 ;
        RECT 11.845 177.435 13.425 177.765 ;
        RECT 20.580 177.435 22.160 177.765 ;
        RECT 29.315 177.435 30.895 177.765 ;
        RECT 38.050 177.435 39.630 177.765 ;
        RECT 27.195 176.050 27.525 176.065 ;
        RECT 27.195 175.750 43.840 176.050 ;
        RECT 27.195 175.735 27.525 175.750 ;
        RECT 15.145 174.715 16.725 175.045 ;
        RECT 23.880 174.715 25.460 175.045 ;
        RECT 32.615 174.715 34.195 175.045 ;
        RECT 41.350 174.715 42.930 175.045 ;
        RECT 43.540 174.690 43.840 175.750 ;
        RECT 44.770 174.690 48.770 174.840 ;
        RECT 43.540 174.390 48.770 174.690 ;
        RECT 44.770 174.240 48.770 174.390 ;
        RECT 46.710 173.140 47.090 173.460 ;
        RECT 2.750 171.290 6.750 171.440 ;
        RECT 18.455 171.290 18.785 171.305 ;
        RECT 2.750 170.990 18.785 171.290 ;
        RECT 2.750 170.840 6.750 170.990 ;
        RECT 18.455 170.975 18.785 170.990 ;
        RECT 46.750 169.965 47.050 173.140 ;
        RECT 46.735 169.635 47.065 169.965 ;
        RECT 14.060 167.890 14.440 167.900 ;
        RECT 19.375 167.890 19.705 167.905 ;
        RECT 14.060 167.590 19.705 167.890 ;
        RECT 14.060 167.580 14.440 167.590 ;
        RECT 19.375 167.575 19.705 167.590 ;
        RECT 23.515 167.890 23.845 167.905 ;
        RECT 44.770 167.890 48.770 168.040 ;
        RECT 23.515 167.590 48.770 167.890 ;
        RECT 23.515 167.575 23.845 167.590 ;
        RECT 44.770 167.440 48.770 167.590 ;
        RECT 27.335 165.950 27.665 165.965 ;
        RECT 1.950 165.650 27.665 165.950 ;
        RECT 27.335 165.635 27.665 165.650 ;
        RECT 47.750 164.670 48.150 164.695 ;
        RECT 46.480 164.320 48.150 164.670 ;
        RECT 47.750 164.295 48.150 164.320 ;
        RECT 48.145 162.475 48.475 162.490 ;
        RECT 49.575 162.475 49.925 162.500 ;
        RECT 48.145 162.175 49.925 162.475 ;
        RECT 48.145 162.160 48.475 162.175 ;
        RECT 49.575 162.150 49.925 162.175 ;
        RECT 47.820 160.950 48.200 160.960 ;
        RECT 51.325 160.950 51.645 160.990 ;
        RECT 47.820 160.650 51.645 160.950 ;
        RECT 47.820 160.640 48.200 160.650 ;
        RECT 51.325 160.610 51.645 160.650 ;
        RECT 46.320 133.765 46.695 133.790 ;
        RECT 44.940 133.440 46.695 133.765 ;
        RECT 46.320 133.415 46.695 133.440 ;
        RECT 47.765 127.980 48.085 128.360 ;
        RECT 47.775 127.220 48.075 127.980 ;
        RECT 47.750 126.870 48.100 127.220 ;
        RECT 53.705 121.645 54.170 196.765 ;
        RECT 57.585 191.400 57.915 191.415 ;
        RECT 62.060 191.400 62.380 191.440 ;
        RECT 57.585 191.100 62.380 191.400 ;
        RECT 57.585 191.085 57.915 191.100 ;
        RECT 62.060 191.060 62.380 191.100 ;
        RECT 63.000 187.700 94.860 196.765 ;
        RECT 62.075 187.540 94.860 187.700 ;
        RECT 62.060 187.200 94.860 187.540 ;
        RECT 62.060 187.190 62.410 187.200 ;
        RECT 63.000 185.000 94.860 187.200 ;
        RECT 96.060 185.000 127.920 213.400 ;
        RECT 129.120 185.000 160.980 213.400 ;
        RECT 54.845 183.260 55.225 183.265 ;
        RECT 56.840 183.260 57.200 183.285 ;
        RECT 54.845 182.950 57.200 183.260 ;
        RECT 54.845 182.945 55.225 182.950 ;
        RECT 56.840 182.925 57.200 182.950 ;
        RECT 63.000 168.635 94.860 183.400 ;
        RECT 40.810 121.180 54.170 121.645 ;
        RECT 54.875 168.170 94.860 168.635 ;
        RECT 54.875 119.985 55.340 168.170 ;
        RECT 58.735 162.535 59.065 162.550 ;
        RECT 61.245 162.535 61.565 162.575 ;
        RECT 58.735 162.235 61.565 162.535 ;
        RECT 58.735 162.220 59.065 162.235 ;
        RECT 61.245 162.195 61.565 162.235 ;
        RECT 55.995 160.950 56.375 160.960 ;
        RECT 57.200 160.950 57.550 160.975 ;
        RECT 55.995 160.650 57.550 160.950 ;
        RECT 55.995 160.640 56.375 160.650 ;
        RECT 57.200 160.625 57.550 160.650 ;
        RECT 63.000 157.700 94.860 168.170 ;
        RECT 61.370 157.610 61.720 157.635 ;
        RECT 62.740 157.610 94.860 157.700 ;
        RECT 61.370 157.310 94.860 157.610 ;
        RECT 61.370 157.285 61.720 157.310 ;
        RECT 62.740 157.200 94.860 157.310 ;
        RECT 56.715 155.065 57.085 155.090 ;
        RECT 55.910 154.745 57.085 155.065 ;
        RECT 63.000 155.000 94.860 157.200 ;
        RECT 96.060 155.000 127.920 183.400 ;
        RECT 129.120 155.000 160.980 183.400 ;
        RECT 56.715 154.720 57.085 154.745 ;
        RECT 63.000 136.820 94.860 153.400 ;
        RECT 35.805 119.520 55.340 119.985 ;
        RECT 55.965 136.355 94.860 136.820 ;
        RECT 55.965 118.535 56.430 136.355 ;
        RECT 57.930 132.670 58.260 132.685 ;
        RECT 60.425 132.670 60.745 132.710 ;
        RECT 57.930 132.370 60.745 132.670 ;
        RECT 57.930 132.355 58.260 132.370 ;
        RECT 60.425 132.330 60.745 132.370 ;
        RECT 61.870 127.700 62.170 127.740 ;
        RECT 63.000 127.700 94.860 136.355 ;
        RECT 61.870 127.260 94.860 127.700 ;
        RECT 61.845 127.200 94.860 127.260 ;
        RECT 61.845 126.910 62.195 127.200 ;
        RECT 63.000 125.000 94.860 127.200 ;
        RECT 96.060 125.000 127.920 153.400 ;
        RECT 129.120 125.000 160.980 153.400 ;
        RECT 20.070 118.070 56.430 118.535 ;
        RECT 20.070 105.185 20.535 118.070 ;
        RECT 63.000 106.270 94.860 123.400 ;
        RECT 22.835 105.805 94.860 106.270 ;
        RECT 8.270 102.340 8.705 102.365 ;
        RECT 6.375 101.955 8.705 102.340 ;
        RECT 8.270 101.930 8.705 101.955 ;
        RECT 22.835 95.100 23.300 105.805 ;
        RECT 46.590 105.015 47.105 105.040 ;
        RECT 46.590 104.550 48.065 105.015 ;
        RECT 46.590 104.525 47.105 104.550 ;
        RECT 56.020 101.055 56.350 101.070 ;
        RECT 59.625 101.055 59.945 101.095 ;
        RECT 56.020 100.755 59.945 101.055 ;
        RECT 56.020 100.740 56.350 100.755 ;
        RECT 59.625 100.715 59.945 100.755 ;
        RECT 35.850 99.560 36.245 99.955 ;
        RECT 38.495 99.855 38.845 99.880 ;
        RECT 39.260 99.855 39.640 99.865 ;
        RECT 35.875 99.100 36.220 99.560 ;
        RECT 38.495 99.555 39.640 99.855 ;
        RECT 40.865 99.735 41.260 100.130 ;
        RECT 43.250 99.895 43.600 99.920 ;
        RECT 44.155 99.895 44.535 99.905 ;
        RECT 38.495 99.530 38.845 99.555 ;
        RECT 39.260 99.545 39.640 99.555 ;
        RECT 40.890 99.100 41.235 99.735 ;
        RECT 43.250 99.595 44.535 99.895 ;
        RECT 45.855 99.810 46.250 100.205 ;
        RECT 43.250 99.570 43.600 99.595 ;
        RECT 44.155 99.585 44.535 99.595 ;
        RECT 45.880 99.100 46.225 99.810 ;
        RECT 20.100 94.635 23.300 95.100 ;
        RECT 27.690 93.780 28.040 93.805 ;
        RECT 30.060 93.780 47.920 99.100 ;
        RECT 53.170 98.020 53.520 98.045 ;
        RECT 27.690 93.480 47.920 93.780 ;
        RECT 51.865 97.720 53.520 98.020 ;
        RECT 51.865 93.640 52.165 97.720 ;
        RECT 53.170 97.695 53.520 97.720 ;
        RECT 63.000 97.700 94.860 105.805 ;
        RECT 62.740 97.605 94.860 97.700 ;
        RECT 61.710 97.255 94.860 97.605 ;
        RECT 62.740 97.200 94.860 97.255 ;
        RECT 53.160 95.305 53.540 95.315 ;
        RECT 54.600 95.305 54.950 95.330 ;
        RECT 53.160 95.005 54.950 95.305 ;
        RECT 53.160 94.995 53.540 95.005 ;
        RECT 54.600 94.980 54.950 95.005 ;
        RECT 63.000 95.000 94.860 97.200 ;
        RECT 96.060 95.000 127.920 123.400 ;
        RECT 129.120 95.000 160.980 123.400 ;
        RECT 27.690 93.455 28.040 93.480 ;
        RECT 6.435 91.220 6.815 91.230 ;
        RECT 8.340 91.220 8.690 91.245 ;
        RECT 6.435 90.920 8.690 91.220 ;
        RECT 6.435 90.910 6.815 90.920 ;
        RECT 8.340 90.895 8.690 90.920 ;
        RECT 27.515 89.580 27.865 89.605 ;
        RECT 30.060 89.580 47.920 93.480 ;
        RECT 51.855 93.260 52.175 93.640 ;
        RECT 27.515 89.280 47.920 89.580 ;
        RECT 27.515 89.255 27.865 89.280 ;
        RECT 27.675 84.975 28.025 85.000 ;
        RECT 30.060 84.975 47.920 89.280 ;
        RECT 27.675 84.675 47.920 84.975 ;
        RECT 27.675 84.650 28.025 84.675 ;
        RECT 30.060 82.700 47.920 84.675 ;
        RECT 33.795 81.735 34.095 82.700 ;
        RECT 37.615 81.805 37.915 82.700 ;
        RECT 33.770 81.385 34.120 81.735 ;
        RECT 35.625 81.360 35.975 81.710 ;
        RECT 37.590 81.455 37.940 81.805 ;
        RECT 41.520 81.430 41.870 81.780 ;
        RECT 44.610 81.740 44.910 82.700 ;
        RECT 35.650 80.980 35.950 81.360 ;
        RECT 41.545 81.015 41.845 81.430 ;
        RECT 44.585 81.390 44.935 81.740 ;
        RECT 35.640 80.600 35.960 80.980 ;
        RECT 41.535 80.635 41.855 81.015 ;
        RECT 6.675 80.080 7.055 80.090 ;
        RECT 8.435 80.080 8.785 80.105 ;
        RECT 6.675 79.780 8.785 80.080 ;
        RECT 6.675 79.770 7.055 79.780 ;
        RECT 8.435 79.755 8.785 79.780 ;
        RECT 45.690 77.170 46.050 77.195 ;
        RECT 46.795 77.170 47.175 77.175 ;
        RECT 45.690 76.860 47.175 77.170 ;
        RECT 45.690 76.835 46.050 76.860 ;
        RECT 46.795 76.855 47.175 76.860 ;
        RECT 63.000 76.000 94.860 93.400 ;
        RECT 20.175 75.535 94.860 76.000 ;
        RECT 4.325 67.805 4.705 67.815 ;
        RECT 25.120 67.805 25.470 67.830 ;
        RECT 4.325 67.505 25.470 67.805 ;
        RECT 4.325 67.495 4.705 67.505 ;
        RECT 25.120 67.480 25.470 67.505 ;
        RECT 30.065 43.740 30.530 74.415 ;
        RECT 45.605 71.990 47.095 72.015 ;
        RECT 45.600 70.490 53.475 71.990 ;
        RECT 55.845 71.535 56.175 71.550 ;
        RECT 58.690 71.535 59.010 71.575 ;
        RECT 55.845 71.235 59.010 71.535 ;
        RECT 55.845 71.220 56.175 71.235 ;
        RECT 58.690 71.195 59.010 71.235 ;
        RECT 45.605 70.465 47.095 70.490 ;
        RECT 52.655 69.165 52.975 69.545 ;
        RECT 52.660 68.295 52.965 69.165 ;
        RECT 52.635 67.940 52.990 68.295 ;
        RECT 63.000 67.700 94.860 75.535 ;
        RECT 62.685 67.695 94.860 67.700 ;
        RECT 61.780 67.270 94.860 67.695 ;
        RECT 62.685 67.200 94.860 67.270 ;
        RECT 52.370 65.590 52.750 65.600 ;
        RECT 54.195 65.590 54.545 65.615 ;
        RECT 52.370 65.290 54.545 65.590 ;
        RECT 52.370 65.280 52.750 65.290 ;
        RECT 54.195 65.265 54.545 65.290 ;
        RECT 63.000 65.000 94.860 67.200 ;
        RECT 96.060 65.000 127.920 93.400 ;
        RECT 129.120 65.000 160.980 93.400 ;
        RECT 63.000 43.740 94.860 63.400 ;
        RECT 30.065 43.275 94.860 43.740 ;
        RECT 55.900 41.885 56.230 41.900 ;
        RECT 57.850 41.885 58.170 41.925 ;
        RECT 55.900 41.585 58.170 41.885 ;
        RECT 55.900 41.570 56.230 41.585 ;
        RECT 57.850 41.545 58.170 41.585 ;
        RECT 38.125 19.040 38.590 41.315 ;
        RECT 53.395 38.795 53.770 38.820 ;
        RECT 47.995 38.470 53.770 38.795 ;
        RECT 53.395 38.445 53.770 38.470 ;
        RECT 63.000 37.700 94.860 43.275 ;
        RECT 61.745 37.200 94.860 37.700 ;
        RECT 52.510 36.075 52.890 36.085 ;
        RECT 54.340 36.075 54.695 36.100 ;
        RECT 52.510 35.770 54.695 36.075 ;
        RECT 52.510 35.765 52.890 35.770 ;
        RECT 54.340 35.745 54.695 35.770 ;
        RECT 63.000 35.000 94.860 37.200 ;
        RECT 96.060 35.000 127.920 63.400 ;
        RECT 129.120 35.000 160.980 63.400 ;
        RECT 63.000 19.040 94.860 33.400 ;
        RECT 38.125 18.575 94.860 19.040 ;
        RECT 56.835 7.850 57.215 8.170 ;
        RECT 56.875 7.215 57.175 7.850 ;
        RECT 63.000 7.700 94.860 18.575 ;
        RECT 46.645 7.080 46.965 7.120 ;
        RECT 54.575 7.080 54.925 7.105 ;
        RECT 46.645 6.780 54.925 7.080 ;
        RECT 56.860 6.885 57.190 7.215 ;
        RECT 61.895 7.200 94.860 7.700 ;
        RECT 46.645 6.740 46.965 6.780 ;
        RECT 54.575 6.755 54.925 6.780 ;
        RECT 61.980 6.625 62.310 7.200 ;
        RECT 63.000 5.000 94.860 7.200 ;
        RECT 96.060 5.000 127.920 33.400 ;
        RECT 129.120 5.000 160.980 33.400 ;
        RECT 54.615 4.300 54.995 4.310 ;
        RECT 55.705 4.300 56.055 4.325 ;
        RECT 54.615 4.000 56.055 4.300 ;
        RECT 54.615 3.990 54.995 4.000 ;
        RECT 55.705 3.975 56.055 4.000 ;
        RECT 152.550 4.145 157.310 4.150 ;
        RECT 152.550 3.255 157.335 4.145 ;
        RECT 152.550 3.250 157.310 3.255 ;
      LAYER met4 ;
        RECT 150.865 224.760 151.190 225.435 ;
        RECT 154.865 224.760 154.870 224.995 ;
        RECT 3.990 223.865 4.290 224.760 ;
        RECT 7.670 223.865 7.970 224.760 ;
        RECT 11.350 223.865 11.650 224.760 ;
        RECT 15.030 223.865 15.330 224.760 ;
        RECT 18.710 223.865 19.010 224.760 ;
        RECT 22.390 223.865 22.690 224.760 ;
        RECT 26.070 223.865 26.370 224.760 ;
        RECT 29.750 223.865 30.050 224.760 ;
        RECT 3.990 223.565 30.050 223.865 ;
        RECT 3.990 220.250 4.290 223.565 ;
        RECT 4.935 222.950 5.265 222.965 ;
        RECT 33.430 222.950 33.730 224.760 ;
        RECT 4.935 222.650 33.730 222.950 ;
        RECT 4.935 222.635 5.265 222.650 ;
        RECT 37.110 222.150 37.410 224.760 ;
        RECT 40.790 223.765 41.090 224.760 ;
        RECT 40.775 223.435 41.105 223.765 ;
        RECT 2.500 219.950 4.290 220.250 ;
        RECT 4.950 221.850 37.410 222.150 ;
        RECT 4.950 200.065 5.250 221.850 ;
        RECT 40.335 220.750 40.665 220.765 ;
        RECT 44.470 220.750 44.770 224.760 ;
        RECT 40.335 220.450 44.770 220.750 ;
        RECT 40.335 220.435 40.665 220.450 ;
        RECT 48.150 219.450 48.450 224.760 ;
        RECT 51.830 223.865 52.130 224.760 ;
        RECT 55.510 223.965 55.810 224.760 ;
        RECT 59.190 223.965 59.490 224.760 ;
        RECT 62.870 224.065 63.170 224.760 ;
        RECT 66.550 224.065 66.850 224.760 ;
        RECT 70.230 224.065 70.530 224.760 ;
        RECT 51.815 223.535 52.145 223.865 ;
        RECT 55.495 223.635 55.825 223.965 ;
        RECT 59.175 223.635 59.505 223.965 ;
        RECT 62.855 223.735 63.185 224.065 ;
        RECT 66.535 223.735 66.865 224.065 ;
        RECT 70.215 223.735 70.545 224.065 ;
        RECT 73.910 223.965 74.210 224.760 ;
        RECT 77.590 224.065 77.890 224.760 ;
        RECT 73.895 223.635 74.225 223.965 ;
        RECT 77.575 223.735 77.905 224.065 ;
        RECT 81.270 223.865 81.570 224.760 ;
        RECT 84.950 223.965 85.250 224.760 ;
        RECT 81.255 223.535 81.585 223.865 ;
        RECT 84.935 223.635 85.265 223.965 ;
        RECT 88.630 221.000 88.930 224.760 ;
        RECT 121.750 224.070 122.050 224.760 ;
        RECT 121.735 223.740 122.065 224.070 ;
        RECT 49.000 220.760 111.465 221.000 ;
        RECT 6.150 219.150 48.450 219.450 ;
        RECT 50.500 219.265 111.465 220.760 ;
        RECT 112.000 220.420 112.330 220.435 ;
        RECT 125.430 220.420 125.730 224.760 ;
        RECT 112.000 220.120 125.730 220.420 ;
        RECT 112.000 220.105 112.330 220.120 ;
        RECT 112.060 219.620 112.390 219.635 ;
        RECT 129.110 219.620 129.410 224.760 ;
        RECT 112.060 219.320 129.410 219.620 ;
        RECT 112.060 219.305 112.390 219.320 ;
        RECT 6.150 208.665 6.450 219.150 ;
        RECT 50.500 218.000 50.610 219.265 ;
        RECT 106.385 218.450 106.715 218.780 ;
        RECT 106.400 217.355 106.700 218.450 ;
        RECT 107.215 217.400 107.545 217.730 ;
        RECT 46.735 216.735 47.065 217.065 ;
        RECT 59.635 217.055 106.700 217.355 ;
        RECT 6.135 208.335 6.465 208.665 ;
        RECT 4.935 199.735 5.265 200.065 ;
        RECT 11.835 175.500 13.435 207.760 ;
        RECT 14.085 195.455 14.415 195.785 ;
        RECT 11.835 174.640 13.500 175.500 ;
        RECT 12.000 174.000 13.500 174.640 ;
        RECT 2.500 172.500 13.500 174.000 ;
        RECT 14.100 167.905 14.400 195.455 ;
        RECT 15.135 174.640 16.735 207.760 ;
        RECT 17.765 189.335 18.095 189.665 ;
        RECT 17.780 178.785 18.080 189.335 ;
        RECT 17.765 178.455 18.095 178.785 ;
        RECT 20.570 174.640 22.170 207.760 ;
        RECT 23.870 174.640 25.470 207.760 ;
        RECT 29.305 174.640 30.905 207.760 ;
        RECT 32.605 174.640 34.205 207.760 ;
        RECT 38.040 174.640 39.640 207.760 ;
        RECT 41.340 174.640 42.940 207.760 ;
        RECT 41.465 172.525 42.850 174.640 ;
        RECT 46.750 173.465 47.050 216.735 ;
        RECT 57.845 216.110 58.175 216.440 ;
        RECT 56.860 211.885 57.190 212.215 ;
        RECT 54.870 183.260 55.200 183.270 ;
        RECT 50.500 182.950 55.200 183.260 ;
        RECT 54.870 182.940 55.200 182.950 ;
        RECT 46.735 173.135 47.065 173.465 ;
        RECT 41.465 170.935 49.000 172.525 ;
        RECT 14.085 167.575 14.415 167.905 ;
        RECT 45.710 160.950 47.210 169.135 ;
        RECT 47.845 160.950 48.175 160.965 ;
        RECT 45.710 160.650 48.175 160.950 ;
        RECT 44.965 133.765 45.300 133.770 ;
        RECT 45.710 133.765 47.210 160.650 ;
        RECT 47.845 160.635 48.175 160.650 ;
        RECT 51.320 160.950 51.650 160.965 ;
        RECT 56.020 160.950 56.350 160.965 ;
        RECT 51.320 160.650 56.350 160.950 ;
        RECT 51.320 160.635 51.650 160.650 ;
        RECT 56.020 160.635 56.350 160.650 ;
        RECT 55.935 155.065 56.265 155.070 ;
        RECT 50.500 154.745 56.265 155.065 ;
        RECT 55.935 154.740 56.265 154.745 ;
        RECT 44.965 133.440 47.210 133.765 ;
        RECT 44.965 133.435 45.300 133.440 ;
        RECT 45.710 130.965 47.210 133.440 ;
        RECT 2.500 129.465 47.210 130.965 ;
        RECT 47.760 128.320 48.090 128.335 ;
        RECT 47.760 128.020 49.000 128.320 ;
        RECT 47.760 128.005 48.090 128.020 ;
        RECT 6.400 102.340 6.795 102.345 ;
        RECT 2.500 101.955 6.795 102.340 ;
        RECT 6.400 101.950 6.795 101.955 ;
        RECT 6.460 91.220 6.790 91.235 ;
        RECT 2.500 90.920 6.790 91.220 ;
        RECT 6.460 90.905 6.790 90.920 ;
        RECT 22.790 83.975 23.635 105.790 ;
        RECT 47.565 105.015 48.040 105.020 ;
        RECT 47.565 104.550 49.000 105.015 ;
        RECT 47.565 104.545 48.040 104.550 ;
        RECT 34.620 100.285 49.000 100.975 ;
        RECT 39.300 99.870 39.600 100.285 ;
        RECT 44.195 99.910 44.495 100.285 ;
        RECT 39.285 99.540 39.615 99.870 ;
        RECT 44.180 99.580 44.510 99.910 ;
        RECT 2.500 83.130 28.075 83.975 ;
        RECT 27.230 81.175 28.075 83.130 ;
        RECT 30.080 82.760 30.560 99.040 ;
        RECT 31.915 92.040 47.525 98.705 ;
        RECT 53.185 95.305 53.515 95.320 ;
        RECT 50.500 95.005 53.515 95.305 ;
        RECT 53.185 94.990 53.515 95.005 ;
        RECT 51.850 93.285 52.180 93.615 ;
        RECT 51.865 92.110 52.165 93.285 ;
        RECT 31.915 90.540 49.000 92.040 ;
        RECT 51.865 91.080 53.445 92.110 ;
        RECT 31.915 83.095 47.525 90.540 ;
        RECT 27.230 80.330 47.125 81.175 ;
        RECT 6.700 80.080 7.030 80.095 ;
        RECT 2.500 79.780 7.030 80.080 ;
        RECT 6.700 79.765 7.030 79.780 ;
        RECT 46.820 77.170 47.150 77.180 ;
        RECT 46.820 76.860 49.000 77.170 ;
        RECT 46.820 76.850 47.150 76.860 ;
        RECT 51.945 71.995 53.445 91.080 ;
        RECT 4.350 67.805 4.680 67.820 ;
        RECT 2.500 67.505 4.680 67.805 ;
        RECT 4.350 67.490 4.680 67.505 ;
        RECT 45.600 38.795 47.100 71.990 ;
        RECT 51.940 70.485 53.450 71.995 ;
        RECT 52.665 69.520 52.970 70.485 ;
        RECT 52.650 69.190 52.980 69.520 ;
        RECT 52.395 65.590 52.725 65.605 ;
        RECT 50.500 65.290 52.725 65.590 ;
        RECT 52.395 65.275 52.725 65.290 ;
        RECT 48.020 38.795 48.355 38.800 ;
        RECT 45.600 38.470 48.355 38.795 ;
        RECT 45.600 10.325 47.100 38.470 ;
        RECT 48.020 38.465 48.355 38.470 ;
        RECT 52.535 36.080 52.865 36.090 ;
        RECT 50.500 35.775 52.865 36.080 ;
        RECT 52.535 35.760 52.865 35.775 ;
        RECT 2.500 8.825 47.100 10.325 ;
        RECT 46.655 7.095 46.955 8.825 ;
        RECT 56.875 8.175 57.175 211.885 ;
        RECT 57.860 41.900 58.160 216.110 ;
        RECT 58.685 215.045 59.015 215.375 ;
        RECT 58.700 71.550 59.000 215.045 ;
        RECT 59.635 101.070 59.935 217.055 ;
        RECT 107.230 216.395 107.530 217.400 ;
        RECT 60.435 216.095 107.530 216.395 ;
        RECT 108.100 216.130 108.430 216.460 ;
        RECT 60.435 132.835 60.735 216.095 ;
        RECT 108.115 215.355 108.415 216.130 ;
        RECT 61.255 215.055 108.415 215.355 ;
        RECT 61.255 162.550 61.555 215.055 ;
        RECT 109.005 214.980 109.335 215.310 ;
        RECT 109.020 214.390 109.320 214.980 ;
        RECT 62.055 214.090 109.320 214.390 ;
        RECT 62.055 213.765 62.715 214.090 ;
        RECT 62.055 213.760 62.370 213.765 ;
        RECT 62.070 191.415 62.370 213.760 ;
        RECT 62.055 191.085 62.385 191.415 ;
        RECT 63.395 185.395 93.005 213.005 ;
        RECT 78.250 183.005 79.750 185.395 ;
        RECT 94.360 185.060 94.840 213.340 ;
        RECT 109.730 213.005 111.465 219.265 ;
        RECT 112.020 218.765 112.350 218.780 ;
        RECT 132.790 218.765 133.090 224.760 ;
        RECT 112.020 218.465 133.090 218.765 ;
        RECT 112.020 218.450 112.350 218.465 ;
        RECT 111.955 217.715 112.285 217.730 ;
        RECT 136.470 217.715 136.770 224.760 ;
        RECT 111.955 217.415 136.770 217.715 ;
        RECT 111.955 217.400 112.285 217.415 ;
        RECT 111.930 216.445 112.260 216.460 ;
        RECT 140.150 216.445 140.450 224.760 ;
        RECT 111.930 216.145 140.450 216.445 ;
        RECT 111.930 216.130 112.260 216.145 ;
        RECT 111.960 215.295 112.290 215.310 ;
        RECT 143.830 215.295 144.130 224.760 ;
        RECT 150.865 215.295 151.485 224.760 ;
        RECT 154.865 222.025 155.165 224.760 ;
        RECT 154.850 221.695 155.180 222.025 ;
        RECT 111.960 214.995 144.130 215.295 ;
        RECT 111.960 214.980 112.290 214.995 ;
        RECT 150.935 214.505 151.420 215.295 ;
        RECT 112.015 214.020 151.420 214.505 ;
        RECT 96.455 185.395 126.065 213.005 ;
        RECT 61.240 162.220 61.570 162.550 ;
        RECT 63.395 155.395 93.005 183.005 ;
        RECT 78.250 153.005 79.750 155.395 ;
        RECT 94.360 155.060 94.840 183.340 ;
        RECT 109.730 183.005 111.465 185.395 ;
        RECT 127.420 185.060 127.900 213.340 ;
        RECT 129.515 185.395 159.125 213.005 ;
        RECT 96.455 155.395 126.065 183.005 ;
        RECT 60.350 132.315 60.810 132.835 ;
        RECT 63.395 125.395 93.005 153.005 ;
        RECT 78.250 123.005 79.750 125.395 ;
        RECT 94.360 125.060 94.840 153.340 ;
        RECT 109.730 153.005 111.465 155.395 ;
        RECT 127.420 155.060 127.900 183.340 ;
        RECT 144.285 183.005 145.785 185.395 ;
        RECT 160.480 185.060 160.960 213.340 ;
        RECT 129.515 155.395 159.125 183.005 ;
        RECT 96.455 125.395 126.065 153.005 ;
        RECT 59.620 100.740 59.950 101.070 ;
        RECT 63.395 95.395 93.005 123.005 ;
        RECT 78.250 93.005 79.750 95.395 ;
        RECT 94.360 95.060 94.840 123.340 ;
        RECT 109.730 123.005 111.465 125.395 ;
        RECT 127.420 125.060 127.900 153.340 ;
        RECT 144.285 153.005 145.785 155.395 ;
        RECT 160.480 155.060 160.960 183.340 ;
        RECT 129.515 125.395 159.125 153.005 ;
        RECT 96.455 95.395 126.065 123.005 ;
        RECT 58.685 71.220 59.015 71.550 ;
        RECT 63.395 65.395 93.005 93.005 ;
        RECT 78.250 63.005 79.750 65.395 ;
        RECT 94.360 65.060 94.840 93.340 ;
        RECT 109.730 93.005 111.465 95.395 ;
        RECT 127.420 95.060 127.900 123.340 ;
        RECT 144.285 123.005 145.785 125.395 ;
        RECT 160.480 125.060 160.960 153.340 ;
        RECT 129.515 95.395 159.125 123.005 ;
        RECT 96.455 65.395 126.065 93.005 ;
        RECT 57.845 41.570 58.175 41.900 ;
        RECT 63.395 35.395 93.005 63.005 ;
        RECT 78.250 33.005 79.750 35.395 ;
        RECT 94.360 35.060 94.840 63.340 ;
        RECT 109.730 63.005 111.465 65.395 ;
        RECT 127.420 65.060 127.900 93.340 ;
        RECT 144.285 93.005 145.785 95.395 ;
        RECT 160.480 95.060 160.960 123.340 ;
        RECT 129.515 65.395 159.125 93.005 ;
        RECT 96.455 35.395 126.065 63.005 ;
        RECT 56.860 7.845 57.190 8.175 ;
        RECT 46.640 6.765 46.970 7.095 ;
        RECT 63.395 5.395 93.005 33.005 ;
        RECT 49.000 4.470 50.500 5.000 ;
        RECT 78.250 4.470 79.750 5.395 ;
        RECT 94.360 5.060 94.840 33.340 ;
        RECT 109.730 33.005 111.465 35.395 ;
        RECT 127.420 35.060 127.900 63.340 ;
        RECT 144.285 63.005 145.785 65.395 ;
        RECT 160.480 65.060 160.960 93.340 ;
        RECT 129.515 35.395 159.125 63.005 ;
        RECT 96.455 5.395 126.065 33.005 ;
        RECT 127.420 5.060 127.900 33.340 ;
        RECT 144.285 33.005 145.785 35.395 ;
        RECT 160.480 35.060 160.960 63.340 ;
        RECT 129.515 5.395 159.125 33.005 ;
        RECT 144.285 4.470 145.785 5.395 ;
        RECT 160.480 5.060 160.960 33.340 ;
        RECT 49.000 2.970 145.785 4.470 ;
        RECT 156.410 1.000 157.310 4.150 ;
  END
END tt_um_adia_psu_full_test
END LIBRARY

