magic
tech sky130A
magscale 1 2
timestamp 1717280941
<< locali >>
rect 11946 37591 12067 37626
rect 11872 37340 11961 37374
rect 11710 37281 11792 37317
rect 11946 37050 12089 37085
rect 11705 31697 11826 31732
rect 11631 31446 11720 31480
rect 11469 31387 11551 31423
rect 11705 31156 11848 31191
rect 11672 25731 11793 25766
rect 11598 25480 11687 25514
rect 11436 25421 11518 25457
rect 11672 25190 11815 25225
rect 3894 20410 4015 20445
rect 6815 20294 7033 20305
rect 6815 20260 9366 20294
rect 6815 20257 7033 20260
rect 7717 20225 7751 20260
rect 3820 20159 3909 20193
rect 8668 20218 8702 20260
rect 3658 20100 3740 20136
rect 3894 19869 4037 19904
rect 4318 19568 4352 19696
rect 11764 19559 11885 19594
rect 11690 19308 11779 19342
rect 11528 19249 11610 19285
rect 11764 19018 11907 19053
rect 3924 18196 4045 18231
rect 3850 17945 3939 17979
rect 3688 17886 3770 17922
rect 3924 17655 4067 17690
rect 4345 17337 4379 17482
rect 3914 15970 4035 16005
rect 6951 15946 6985 15977
rect 6285 15912 7329 15946
rect 7766 15898 8066 15932
rect 8100 15898 8696 15932
rect 5652 15828 5788 15863
rect 7162 15817 7298 15852
rect 8561 15817 8697 15852
rect 3840 15719 3929 15753
rect 3678 15660 3760 15696
rect 5576 15577 5665 15615
rect 7086 15566 7175 15604
rect 8485 15566 8574 15604
rect 5435 15524 5499 15561
rect 6945 15513 7009 15550
rect 8344 15513 8408 15550
rect 3914 15429 4057 15464
rect 4338 15234 4439 15268
rect 11664 13606 11785 13641
rect 11590 13355 11679 13389
rect 11428 13296 11510 13332
rect 11664 13065 11807 13100
rect 11638 7707 11759 7742
rect 11564 7456 11653 7490
rect 11402 7397 11484 7433
rect 11638 7166 11781 7201
rect 11844 1364 11965 1399
rect 11770 1113 11859 1147
rect 11608 1054 11690 1090
rect 11844 823 11987 858
<< viali >>
rect 11961 37340 11995 37374
rect 11674 37281 11710 37317
rect 11720 31446 11754 31480
rect 11433 31387 11469 31423
rect 11687 25480 11721 25514
rect 11400 25421 11436 25457
rect 6767 20257 6815 20305
rect 3909 20159 3943 20193
rect 7717 20191 7751 20225
rect 8668 20184 8702 20218
rect 3622 20100 3658 20136
rect 4318 19534 4352 19568
rect 11779 19308 11813 19342
rect 11492 19249 11528 19285
rect 3939 17945 3973 17979
rect 3652 17886 3688 17922
rect 4345 17303 4379 17337
rect 6951 15977 6985 16011
rect 8066 15898 8100 15932
rect 3929 15719 3963 15753
rect 3642 15660 3678 15696
rect 5665 15577 5703 15615
rect 7175 15566 7213 15604
rect 8574 15566 8612 15604
rect 5398 15524 5435 15561
rect 6908 15513 6945 15550
rect 8307 15513 8344 15550
rect 4439 15234 4473 15268
rect 11679 13355 11713 13389
rect 11392 13296 11428 13332
rect 11653 7456 11687 7490
rect 11366 7397 11402 7433
rect 11859 1113 11893 1147
rect 11572 1054 11608 1090
<< metal1 >>
rect 11670 44490 11730 44496
rect 11210 44430 11670 44490
rect 9590 43890 9650 43896
rect 10270 43890 10330 43896
rect 9650 43830 10270 43890
rect 9590 43824 9650 43830
rect 10270 43824 10330 43830
rect 11210 42850 11270 44430
rect 11670 44424 11730 44430
rect 11210 42784 11270 42790
rect 11050 42630 11110 42636
rect 9424 42570 9430 42630
rect 9490 42570 11050 42630
rect 11050 42564 11110 42570
rect 10850 42410 10910 42416
rect 9424 42350 9430 42410
rect 9490 42350 10850 42410
rect 10850 42344 10910 42350
rect 10650 39010 10710 39016
rect 9504 38950 9510 39010
rect 9570 38950 10650 39010
rect 10650 38944 10710 38950
rect 12192 37979 12268 38049
rect 11049 37572 11751 37642
rect 10470 34930 10530 34936
rect 9564 34870 9570 34930
rect 9630 34870 10470 34930
rect 10470 34864 10530 34870
rect 9555 33706 9625 33712
rect 11049 33706 11119 37572
rect 12088 37534 12180 37566
rect 12274 37534 12340 37566
rect 12088 37499 12120 37534
rect 12078 37493 12130 37499
rect 12078 37435 12130 37441
rect 11955 37374 12001 37386
rect 12217 37374 12251 37500
rect 11955 37340 11961 37374
rect 11995 37340 12251 37374
rect 11514 37273 11520 37333
rect 11580 37329 11689 37333
rect 11580 37317 11716 37329
rect 11955 37328 12001 37340
rect 11580 37281 11674 37317
rect 11710 37281 11716 37317
rect 11580 37273 11716 37281
rect 11668 37269 11716 37273
rect 12308 37322 12340 37534
rect 12421 37332 12473 37338
rect 12308 37290 12421 37322
rect 11674 37185 11710 37269
rect 11674 37149 12254 37185
rect 11373 37101 11435 37107
rect 12308 37103 12340 37290
rect 12421 37274 12473 37280
rect 11435 37039 11747 37101
rect 12256 37071 12340 37103
rect 11373 37033 11435 37039
rect 12088 37035 12198 37067
rect 12088 36977 12120 37035
rect 12072 36925 12078 36977
rect 12130 36925 12136 36977
rect 12190 36919 12266 36989
rect 9625 33636 11119 33706
rect 9555 33630 9625 33636
rect 10090 33390 10150 33396
rect 8764 33330 8770 33390
rect 8830 33330 10090 33390
rect 10090 33324 10150 33330
rect 11200 32690 11280 32700
rect 9544 32630 9550 32690
rect 9610 32630 11210 32690
rect 11270 32630 11280 32690
rect 11200 32620 11280 32630
rect 11377 32507 11437 32513
rect 11201 32447 11377 32507
rect 11201 31429 11261 32447
rect 11377 32441 11437 32447
rect 11951 32085 12027 32155
rect 11443 31918 11449 31970
rect 11501 31918 11507 31970
rect 11451 31696 11499 31918
rect 11847 31640 11939 31672
rect 12033 31640 12099 31672
rect 11847 31605 11879 31640
rect 11837 31599 11889 31605
rect 11837 31541 11889 31547
rect 11714 31480 11760 31492
rect 11976 31480 12010 31606
rect 11714 31446 11720 31480
rect 11754 31446 12010 31480
rect 11427 31429 11475 31435
rect 11714 31434 11760 31446
rect 11201 31423 11475 31429
rect 11201 31387 11433 31423
rect 11469 31387 11475 31423
rect 11201 31375 11475 31387
rect 12067 31420 12099 31640
rect 12283 31430 12335 31436
rect 12067 31388 12283 31420
rect 11201 31369 11469 31375
rect 11433 31291 11469 31369
rect 11433 31255 12013 31291
rect 12067 31209 12099 31388
rect 12283 31372 12335 31378
rect 11342 31137 11348 31201
rect 11412 31137 11507 31201
rect 12015 31177 12099 31209
rect 11847 31141 11957 31173
rect 11847 31083 11879 31141
rect 11831 31031 11837 31083
rect 11889 31031 11895 31083
rect 11949 31025 12025 31095
rect 9544 26688 9550 26753
rect 9615 26688 11637 26753
rect 11386 26534 11446 26540
rect 11215 26474 11386 26534
rect 11215 25464 11275 26474
rect 11386 26468 11446 26474
rect 11572 26040 11637 26688
rect 11918 26119 11994 26189
rect 11410 25975 11637 26040
rect 11410 25721 11475 25975
rect 11814 25674 11906 25706
rect 12000 25674 12066 25706
rect 11814 25639 11846 25674
rect 11804 25633 11856 25639
rect 11804 25575 11856 25581
rect 11681 25514 11727 25526
rect 11943 25514 11977 25640
rect 11681 25480 11687 25514
rect 11721 25480 11977 25514
rect 11394 25464 11442 25469
rect 11681 25468 11727 25480
rect 11215 25457 11442 25464
rect 11215 25421 11400 25457
rect 11436 25421 11442 25457
rect 11215 25409 11442 25421
rect 12034 25433 12066 25674
rect 12258 25443 12310 25449
rect 11215 25404 11436 25409
rect 11400 25325 11436 25404
rect 12034 25401 12258 25433
rect 11400 25289 11980 25325
rect 12034 25243 12066 25401
rect 12258 25385 12310 25391
rect 9556 25232 9614 25238
rect 9614 25174 11471 25232
rect 11982 25211 12066 25243
rect 11814 25175 11924 25207
rect 9556 25168 9614 25174
rect 11814 25117 11846 25175
rect 11798 25065 11804 25117
rect 11856 25065 11862 25117
rect 11916 25059 11992 25129
rect 8160 22891 8253 22897
rect 7165 22796 7171 22889
rect 7264 22796 7270 22889
rect 7171 22724 7264 22796
rect 7170 22672 7264 22724
rect 8160 22678 8253 22798
rect 4140 20798 4216 20868
rect 7170 20491 7246 22672
rect 8173 20488 8238 22678
rect 9153 20910 9159 21003
rect 9252 20910 9258 21003
rect 9159 20483 9252 20910
rect 1996 20391 2002 20468
rect 2079 20391 3703 20468
rect 7078 20405 7138 20477
rect 8681 20475 8741 20481
rect 7280 20414 7505 20474
rect 7565 20414 7571 20474
rect 8085 20402 8145 20474
rect 8292 20415 8681 20475
rect 8681 20409 8741 20415
rect 9075 20396 9135 20468
rect 9618 20467 9678 20473
rect 9280 20407 9618 20467
rect 9618 20401 9678 20407
rect 4036 20353 4128 20385
rect 4222 20353 4288 20385
rect 4036 20318 4068 20353
rect 4026 20312 4078 20318
rect 4026 20254 4078 20260
rect 3903 20193 3949 20205
rect 4165 20193 4199 20319
rect 3903 20159 3909 20193
rect 3943 20159 4199 20193
rect 3616 20136 3664 20148
rect 3903 20147 3949 20159
rect 3616 20100 3622 20136
rect 3658 20100 3664 20136
rect 4256 20133 4288 20353
rect 6558 20255 6564 20307
rect 6616 20305 6622 20307
rect 6761 20305 6821 20317
rect 6616 20257 6767 20305
rect 6815 20257 6821 20305
rect 6616 20255 6622 20257
rect 6761 20245 6821 20257
rect 7175 20183 7244 20375
rect 7705 20225 7763 20231
rect 7705 20191 7717 20225
rect 7751 20191 7763 20225
rect 7705 20185 7763 20191
rect 8178 20189 8247 20381
rect 3616 20088 3664 20100
rect 4250 20088 4829 20133
rect 7717 20134 7751 20185
rect 7175 20108 7244 20114
rect 7708 20128 7760 20134
rect 3455 20027 3515 20033
rect 3622 20027 3658 20088
rect 3515 20004 3658 20027
rect 3515 19968 4202 20004
rect 3515 19967 3654 19968
rect 3455 19961 3515 19967
rect 4256 19922 4288 20088
rect 4204 19890 4288 19922
rect 4036 19854 4146 19886
rect 4036 19796 4068 19854
rect 4020 19744 4026 19796
rect 4078 19744 4084 19796
rect 4138 19738 4214 19808
rect 4306 19568 4364 19574
rect 4306 19534 4318 19568
rect 4352 19534 4364 19568
rect 4306 19528 4364 19534
rect 4318 19444 4352 19528
rect 4309 19438 4361 19444
rect 4309 19380 4361 19386
rect 4784 18747 4829 20088
rect 8656 20218 8714 20224
rect 8656 20184 8668 20218
rect 8702 20184 8714 20218
rect 8656 20178 8714 20184
rect 9176 20186 9245 20378
rect 8668 20125 8702 20178
rect 8178 20114 8247 20120
rect 8659 20119 8711 20125
rect 7708 20070 7760 20076
rect 9176 20111 9245 20117
rect 8659 20061 8711 20067
rect 12010 19947 12086 20017
rect 10948 19544 10954 19604
rect 11014 19544 11564 19604
rect 11906 19502 11998 19534
rect 12092 19502 12158 19534
rect 11906 19467 11938 19502
rect 11896 19461 11948 19467
rect 11896 19403 11948 19409
rect 11773 19342 11819 19354
rect 12035 19342 12069 19468
rect 11773 19308 11779 19342
rect 11813 19308 12069 19342
rect 11201 19241 11207 19301
rect 11267 19297 11505 19301
rect 11267 19285 11534 19297
rect 11773 19296 11819 19308
rect 11267 19249 11492 19285
rect 11528 19249 11534 19285
rect 11267 19241 11534 19249
rect 11486 19237 11534 19241
rect 12126 19294 12158 19502
rect 12351 19304 12403 19310
rect 12126 19262 12351 19294
rect 11492 19153 11528 19237
rect 11492 19117 12072 19153
rect 12126 19071 12158 19262
rect 12351 19246 12403 19252
rect 11179 19001 11185 19060
rect 11244 19001 11564 19060
rect 12074 19039 12158 19071
rect 11906 19003 12016 19035
rect 11906 18945 11938 19003
rect 11890 18893 11896 18945
rect 11948 18893 11954 18945
rect 12008 18887 12084 18957
rect 5204 18747 5210 18751
rect 4784 18702 5210 18747
rect 5204 18699 5210 18702
rect 5262 18699 5268 18751
rect 4170 18584 4246 18654
rect 2025 18184 2031 18244
rect 2091 18184 3724 18244
rect 4066 18139 4158 18171
rect 4252 18139 4318 18171
rect 4066 18104 4098 18139
rect 4056 18098 4108 18104
rect 4056 18040 4108 18046
rect 3933 17979 3979 17991
rect 4195 17979 4229 18105
rect 3933 17945 3939 17979
rect 3973 17945 4229 17979
rect 3646 17922 3694 17934
rect 3933 17933 3979 17945
rect 3646 17886 3652 17922
rect 3688 17886 3694 17922
rect 4286 17908 4318 18139
rect 5179 17908 5185 17912
rect 3646 17874 3694 17886
rect 3229 17807 3289 17813
rect 3652 17807 3688 17874
rect 4280 17864 5185 17908
rect 3289 17790 3688 17807
rect 3289 17754 4232 17790
rect 3289 17747 3681 17754
rect 3229 17741 3289 17747
rect 4286 17708 4318 17864
rect 5179 17860 5185 17864
rect 5237 17860 5243 17912
rect 4234 17676 4318 17708
rect 4066 17640 4176 17672
rect 4066 17582 4098 17640
rect 4050 17530 4056 17582
rect 4108 17530 4114 17582
rect 4168 17524 4244 17594
rect 4333 17337 4391 17343
rect 4333 17303 4345 17337
rect 4379 17303 4391 17337
rect 4333 17297 4391 17303
rect 4345 17219 4379 17297
rect 4336 17213 4388 17219
rect 4336 17155 4388 17161
rect 5197 16985 5203 16990
rect 4823 16942 5203 16985
rect 4160 16358 4236 16428
rect 1967 15959 1973 16013
rect 2027 15959 3711 16013
rect 4056 15913 4148 15945
rect 4242 15913 4308 15945
rect 4056 15878 4088 15913
rect 4046 15872 4098 15878
rect 4046 15814 4098 15820
rect 3923 15753 3969 15765
rect 4185 15753 4219 15879
rect 3923 15719 3929 15753
rect 3963 15719 4219 15753
rect 3636 15696 3684 15708
rect 3923 15707 3969 15719
rect 4276 15701 4308 15913
rect 4823 15701 4866 16942
rect 5197 16938 5203 16942
rect 5255 16938 5261 16990
rect 6942 16333 6994 16339
rect 8051 16295 8057 16347
rect 8109 16295 8115 16347
rect 6942 16275 6994 16281
rect 6013 16063 6759 16122
rect 6818 16063 6824 16122
rect 6013 15804 6072 16063
rect 6951 16017 6985 16275
rect 7523 16094 7582 16100
rect 6939 16011 6997 16017
rect 6939 15977 6951 16011
rect 6985 15977 6997 16011
rect 6939 15971 6997 15977
rect 3636 15660 3642 15696
rect 3678 15660 3684 15696
rect 3636 15648 3684 15660
rect 4271 15658 4866 15701
rect 3022 15587 3082 15593
rect 3642 15587 3678 15648
rect 3082 15564 3678 15587
rect 3082 15528 4222 15564
rect 3082 15527 3669 15528
rect 3022 15521 3082 15527
rect 4276 15482 4308 15658
rect 5659 15615 5709 15627
rect 5852 15615 5890 15792
rect 6178 15739 6234 15803
rect 7523 15793 7582 16035
rect 8066 15938 8100 16295
rect 8922 16113 8981 16119
rect 8054 15932 8112 15938
rect 8054 15898 8066 15932
rect 8100 15898 8112 15932
rect 8054 15892 8112 15898
rect 8922 15793 8981 16054
rect 5055 15575 5115 15581
rect 5659 15577 5665 15615
rect 5703 15577 5890 15615
rect 5115 15564 5356 15575
rect 5392 15564 5441 15573
rect 5659 15565 5709 15577
rect 5115 15561 5441 15564
rect 5115 15524 5398 15561
rect 5435 15524 5441 15561
rect 5115 15521 5441 15524
rect 5115 15515 5356 15521
rect 5055 15509 5115 15515
rect 5392 15512 5441 15521
rect 6015 15519 6074 15735
rect 7169 15604 7219 15616
rect 7362 15604 7400 15781
rect 7688 15728 7744 15792
rect 7169 15566 7175 15604
rect 7213 15566 7400 15604
rect 6607 15558 6667 15564
rect 4224 15450 4308 15482
rect 4056 15414 4166 15446
rect 4056 15356 4088 15414
rect 4040 15304 4046 15356
rect 4098 15304 4104 15356
rect 4158 15298 4234 15368
rect 4602 15358 4654 15364
rect 6013 15349 6106 15519
rect 6667 15553 6854 15558
rect 6902 15553 6951 15562
rect 7169 15554 7219 15566
rect 6667 15550 6951 15553
rect 6667 15513 6908 15550
rect 6945 15513 6951 15550
rect 7525 15514 7584 15724
rect 8568 15604 8618 15616
rect 8761 15604 8799 15781
rect 9087 15728 9143 15792
rect 8924 15611 8983 15724
rect 8568 15566 8574 15604
rect 8612 15566 8799 15604
rect 8060 15548 8120 15554
rect 8301 15553 8350 15562
rect 8568 15554 8618 15566
rect 8222 15550 8350 15553
rect 8925 15552 8983 15611
rect 8222 15548 8307 15550
rect 6667 15510 6951 15513
rect 6667 15498 6854 15510
rect 6902 15501 6951 15510
rect 6607 15492 6667 15498
rect 7517 15383 7610 15514
rect 8120 15513 8307 15548
rect 8344 15513 8350 15550
rect 8120 15510 8350 15513
rect 8120 15488 8252 15510
rect 8301 15501 8350 15510
rect 8924 15494 8983 15552
rect 8060 15482 8120 15488
rect 4602 15300 4654 15306
rect 4433 15268 4479 15280
rect 4611 15268 4645 15300
rect 4433 15234 4439 15268
rect 4473 15234 4645 15268
rect 4433 15222 4479 15234
rect 5611 15009 5673 15302
rect 6007 15256 6013 15349
rect 6106 15256 6112 15349
rect 6927 15256 7178 15318
rect 7517 15290 7718 15383
rect 6927 15009 6989 15256
rect 5611 14947 6989 15009
rect 7116 13716 7178 15256
rect 7625 13941 7718 15290
rect 8321 15256 8676 15318
rect 8738 15256 8744 15318
rect 7619 13848 7625 13941
rect 7718 13848 7724 13941
rect 8321 13716 8383 15256
rect 7116 13654 8383 13716
rect 8925 13560 8983 15494
rect 11910 13994 11986 14064
rect 10818 13593 10824 13654
rect 10885 13593 11465 13654
rect 5524 13502 5530 13560
rect 5588 13502 8983 13560
rect 11806 13549 11898 13581
rect 11992 13549 12058 13581
rect 11806 13514 11838 13549
rect 11796 13508 11848 13514
rect 11796 13450 11848 13456
rect 11673 13389 11719 13401
rect 11935 13389 11969 13515
rect 11673 13355 11679 13389
rect 11713 13355 11969 13389
rect 11166 13289 11172 13349
rect 11232 13344 11402 13349
rect 11232 13332 11434 13344
rect 11673 13343 11719 13355
rect 11232 13296 11392 13332
rect 11428 13296 11434 13332
rect 11232 13289 11434 13296
rect 11386 13284 11434 13289
rect 12026 13335 12058 13549
rect 12232 13335 12238 13345
rect 12026 13303 12238 13335
rect 11392 13200 11428 13284
rect 11392 13164 11972 13200
rect 12026 13118 12058 13303
rect 12232 13293 12238 13303
rect 12290 13293 12296 13345
rect 11150 13059 11156 13117
rect 11214 13059 11463 13117
rect 11974 13086 12058 13118
rect 11806 13050 11916 13082
rect 11806 12992 11838 13050
rect 11790 12940 11796 12992
rect 11848 12940 11854 12992
rect 11908 12934 11984 13004
rect 11884 8095 11960 8165
rect 10936 7694 10942 7759
rect 11007 7694 11441 7759
rect 11780 7650 11872 7682
rect 11966 7650 12032 7682
rect 11780 7615 11812 7650
rect 11770 7609 11822 7615
rect 11770 7551 11822 7557
rect 11647 7490 11693 7502
rect 11909 7490 11943 7616
rect 11647 7456 11653 7490
rect 11687 7456 11943 7490
rect 11360 7440 11408 7445
rect 11647 7444 11693 7456
rect 11177 7380 11183 7440
rect 11243 7433 11408 7440
rect 11243 7397 11366 7433
rect 11402 7397 11408 7433
rect 11243 7385 11408 7397
rect 12000 7388 12032 7650
rect 12232 7388 12238 7398
rect 11243 7380 11402 7385
rect 11366 7301 11402 7380
rect 12000 7356 12238 7388
rect 11366 7265 11946 7301
rect 12000 7219 12032 7356
rect 12232 7346 12238 7356
rect 12290 7346 12296 7398
rect 11176 7154 11182 7215
rect 11243 7154 11439 7215
rect 11948 7187 12032 7219
rect 11780 7151 11890 7183
rect 11780 7093 11812 7151
rect 11764 7041 11770 7093
rect 11822 7041 11828 7093
rect 11882 7035 11958 7105
rect 12090 1752 12166 1822
rect 11171 1356 11177 1415
rect 11236 1356 11644 1415
rect 11986 1307 12078 1339
rect 12172 1307 12238 1339
rect 11986 1272 12018 1307
rect 11976 1266 12028 1272
rect 11976 1208 12028 1214
rect 11853 1147 11899 1159
rect 12115 1147 12149 1273
rect 11853 1113 11859 1147
rect 11893 1113 12149 1147
rect 12206 1150 12238 1307
rect 11369 1051 11375 1111
rect 11435 1102 11601 1111
rect 11435 1090 11614 1102
rect 11853 1101 11899 1113
rect 11435 1054 11572 1090
rect 11608 1054 11614 1090
rect 11435 1051 11614 1054
rect 11566 1042 11614 1051
rect 12206 1084 12396 1150
rect 12462 1084 12468 1150
rect 11572 958 11608 1042
rect 11572 922 12152 958
rect 12206 876 12238 1084
rect 11361 800 11367 860
rect 11427 800 11644 860
rect 12154 844 12238 876
rect 11986 808 12096 840
rect 11986 750 12018 808
rect 11970 698 11976 750
rect 12028 698 12034 750
rect 12088 692 12164 762
<< via1 >>
rect 11670 44430 11730 44490
rect 9590 43830 9650 43890
rect 10270 43830 10330 43890
rect 11210 42790 11270 42850
rect 9430 42570 9490 42630
rect 11050 42570 11110 42630
rect 9430 42350 9490 42410
rect 10850 42350 10910 42410
rect 9510 38950 9570 39010
rect 10650 38950 10710 39010
rect 9570 34870 9630 34930
rect 10470 34870 10530 34930
rect 12078 37441 12130 37493
rect 11520 37273 11580 37333
rect 12421 37280 12473 37332
rect 11373 37039 11435 37101
rect 12078 36925 12130 36977
rect 9555 33636 9625 33706
rect 8770 33330 8830 33390
rect 10090 33330 10150 33390
rect 9550 32630 9610 32690
rect 11210 32630 11270 32690
rect 11377 32447 11437 32507
rect 11449 31918 11501 31970
rect 11837 31547 11889 31599
rect 12283 31378 12335 31430
rect 11348 31137 11412 31201
rect 11837 31031 11889 31083
rect 9550 26688 9615 26753
rect 11386 26474 11446 26534
rect 11804 25581 11856 25633
rect 12258 25391 12310 25443
rect 9556 25174 9614 25232
rect 11804 25065 11856 25117
rect 7171 22796 7264 22889
rect 8160 22798 8253 22891
rect 9159 20910 9252 21003
rect 2002 20391 2079 20468
rect 7505 20414 7565 20474
rect 8681 20415 8741 20475
rect 9618 20407 9678 20467
rect 4026 20260 4078 20312
rect 6564 20255 6616 20307
rect 7175 20114 7244 20183
rect 3455 19967 3515 20027
rect 4026 19744 4078 19796
rect 4309 19386 4361 19438
rect 7708 20076 7760 20128
rect 8178 20120 8247 20189
rect 8659 20067 8711 20119
rect 9176 20117 9245 20186
rect 10954 19544 11014 19604
rect 11896 19409 11948 19461
rect 11207 19241 11267 19301
rect 12351 19252 12403 19304
rect 11185 19001 11244 19060
rect 11896 18893 11948 18945
rect 5210 18699 5262 18751
rect 2031 18184 2091 18244
rect 4056 18046 4108 18098
rect 3229 17747 3289 17807
rect 5185 17860 5237 17912
rect 4056 17530 4108 17582
rect 4336 17161 4388 17213
rect 1973 15959 2027 16013
rect 4046 15820 4098 15872
rect 5203 16938 5255 16990
rect 6942 16281 6994 16333
rect 8057 16295 8109 16347
rect 6759 16063 6818 16122
rect 7523 16035 7582 16094
rect 3022 15527 3082 15587
rect 8922 16054 8981 16113
rect 5055 15515 5115 15575
rect 4046 15304 4098 15356
rect 4602 15306 4654 15358
rect 6607 15498 6667 15558
rect 8060 15488 8120 15548
rect 6013 15256 6106 15349
rect 8676 15256 8738 15318
rect 7625 13848 7718 13941
rect 10824 13593 10885 13654
rect 5530 13502 5588 13560
rect 11796 13456 11848 13508
rect 11172 13289 11232 13349
rect 12238 13293 12290 13345
rect 11156 13059 11214 13117
rect 11796 12940 11848 12992
rect 10942 7694 11007 7759
rect 11770 7557 11822 7609
rect 11183 7380 11243 7440
rect 12238 7346 12290 7398
rect 11182 7154 11243 7215
rect 11770 7041 11822 7093
rect 11177 1356 11236 1415
rect 11976 1214 12028 1266
rect 11375 1051 11435 1111
rect 12396 1084 12462 1150
rect 11367 800 11427 860
rect 11976 698 12028 750
<< metal2 >>
rect 9350 44768 9410 44770
rect 9343 44712 9352 44768
rect 9408 44712 9417 44768
rect 6632 44150 6688 44157
rect 6370 44148 6690 44150
rect 6370 44092 6632 44148
rect 6688 44092 6690 44148
rect 6370 44090 6690 44092
rect 8294 44140 8354 44149
rect 6632 44083 6688 44090
rect 8294 44071 8354 44080
rect 3150 43728 3210 43910
rect 3143 43672 3152 43728
rect 3208 43672 3217 43728
rect 3150 43670 3210 43672
rect 9350 43650 9410 44712
rect 24350 44657 24410 44659
rect 12574 44628 12634 44630
rect 14046 44628 14106 44630
rect 14782 44628 14842 44630
rect 11838 44608 11898 44610
rect 9752 44590 9808 44597
rect 9750 44588 9810 44590
rect 9750 44532 9752 44588
rect 9808 44532 9810 44588
rect 11831 44552 11840 44608
rect 11896 44552 11905 44608
rect 12567 44572 12576 44628
rect 12632 44572 12641 44628
rect 13310 44608 13370 44610
rect 9584 43830 9590 43890
rect 9650 43830 9656 43890
rect 9590 43670 9650 43830
rect 9350 43581 9410 43590
rect 9430 42630 9490 42636
rect 9121 42570 9130 42630
rect 9190 42570 9430 42630
rect 9430 42564 9490 42570
rect 9430 42410 9490 42416
rect 9281 42350 9290 42410
rect 9350 42350 9430 42410
rect 9430 42344 9490 42350
rect 9510 39010 9570 39016
rect 9361 38950 9370 39010
rect 9430 38950 9510 39010
rect 9510 38944 9570 38950
rect 941 37610 950 37670
rect 1010 37610 1019 37670
rect 761 34210 770 34270
rect 830 34210 839 34270
rect 770 32310 830 34210
rect 950 32490 1010 37610
rect 1121 36230 1130 36290
rect 1190 36230 1199 36290
rect 1130 32690 1190 36230
rect 9570 34930 9630 34936
rect 9421 34870 9430 34930
rect 9490 34870 9570 34930
rect 9570 34864 9630 34870
rect 9350 33988 9410 33990
rect 9343 33932 9352 33988
rect 9408 33932 9417 33988
rect 8770 33390 8830 33396
rect 7010 33330 8770 33390
rect 8770 33324 8830 33330
rect 5472 33190 5528 33197
rect 9350 33190 9410 33932
rect 9549 33636 9555 33706
rect 9625 33636 9631 33706
rect 5470 33188 5770 33190
rect 5470 33132 5472 33188
rect 5528 33132 5770 33188
rect 5470 33130 5770 33132
rect 8950 33130 9410 33190
rect 5472 33123 5528 33130
rect 9555 32934 9625 33636
rect 9546 32864 9555 32934
rect 9625 32864 9634 32934
rect 9550 32690 9610 32696
rect 1130 32630 9550 32690
rect 9550 32624 9610 32630
rect 9634 32495 9690 32502
rect 9532 32493 9692 32495
rect 9532 32490 9634 32493
rect 950 32437 9634 32490
rect 9690 32437 9692 32493
rect 9750 32490 9810 44532
rect 11838 44490 11898 44552
rect 11664 44430 11670 44490
rect 11730 44430 11898 44490
rect 12574 44330 12634 44572
rect 13303 44552 13312 44608
rect 13368 44552 13377 44608
rect 14039 44572 14048 44628
rect 14104 44572 14113 44628
rect 14775 44572 14784 44628
rect 14840 44572 14849 44628
rect 15518 44608 15578 44610
rect 16254 44608 16314 44610
rect 9950 44320 12634 44330
rect 9920 44270 12634 44320
rect 9920 32495 9980 44270
rect 13310 44110 13370 44552
rect 10090 44050 13370 44110
rect 10090 33390 10150 44050
rect 14046 43890 14106 44572
rect 10264 43830 10270 43890
rect 10330 43830 14106 43890
rect 10084 33330 10090 33390
rect 10150 33330 10156 33390
rect 950 32435 9692 32437
rect 950 32430 9595 32435
rect 9634 32428 9690 32435
rect 9743 32430 9812 32490
rect 9911 32435 9920 32495
rect 9980 32435 9989 32495
rect 9917 32430 9980 32435
rect 9750 32310 9810 32430
rect 770 32250 9810 32310
rect 9550 26753 9615 26759
rect 9260 26688 9269 26753
rect 9334 26688 9550 26753
rect 9550 26682 9615 26688
rect 9555 25439 9615 25448
rect 9555 25370 9615 25379
rect 9556 25232 9614 25370
rect 9550 25174 9556 25232
rect 9614 25174 9620 25232
rect 8162 24324 8255 24329
rect 8158 24241 8167 24324
rect 8250 24241 8259 24324
rect 7161 23992 7254 23997
rect 7157 23909 7166 23992
rect 7249 23909 7258 23992
rect 7161 23297 7254 23909
rect 8162 23297 8255 24241
rect 7161 23200 7264 23297
rect 7171 22889 7264 23200
rect 8160 23194 8255 23297
rect 8160 22891 8253 23194
rect 8154 22798 8160 22891
rect 8253 22798 8259 22891
rect 7171 22790 7264 22796
rect 9750 22641 9810 32250
rect 2323 22581 9810 22641
rect 2002 20468 2079 20474
rect 1650 20391 1659 20468
rect 1736 20391 2002 20468
rect 2002 20385 2079 20391
rect 2031 18244 2091 18250
rect 1664 18184 1673 18244
rect 1733 18184 2031 18244
rect 2031 18178 2091 18184
rect 1683 15956 1692 16016
rect 1752 16013 1761 16016
rect 1973 16013 2027 16019
rect 1752 15959 1973 16013
rect 1752 15956 1761 15959
rect 1973 15953 2027 15959
rect 2323 14350 2383 22581
rect 9920 22347 9980 32430
rect 2582 22287 9980 22347
rect 2582 14675 2642 22287
rect 10090 22096 10150 33330
rect 2794 22036 10150 22096
rect 2794 14922 2854 22036
rect 10270 21795 10330 43830
rect 14782 43690 14842 44572
rect 15511 44552 15520 44608
rect 15576 44552 15585 44608
rect 16247 44552 16256 44608
rect 16312 44552 16321 44608
rect 24343 44601 24352 44657
rect 24408 44601 24417 44657
rect 16990 44568 17050 44570
rect 10470 43630 14842 43690
rect 10470 34930 10530 43630
rect 15518 43490 15578 44552
rect 10650 43430 15578 43490
rect 10650 39010 10710 43430
rect 16254 43290 16314 44552
rect 16983 44512 16992 44568
rect 17048 44512 17057 44568
rect 10850 43230 16314 43290
rect 10850 42410 10910 43230
rect 16990 43110 17050 44512
rect 11050 43050 17050 43110
rect 11050 42630 11110 43050
rect 24350 42862 24410 44601
rect 11204 42790 11210 42850
rect 11270 42790 11276 42850
rect 11375 42802 24410 42862
rect 11044 42570 11050 42630
rect 11110 42570 11116 42630
rect 10844 42350 10850 42410
rect 10910 42350 10916 42410
rect 10644 38950 10650 39010
rect 10710 38950 10716 39010
rect 10464 34870 10470 34930
rect 10530 34870 10536 34930
rect 3022 21735 10330 21795
rect 3022 15587 3082 21735
rect 10470 21529 10530 34870
rect 3229 21469 10530 21529
rect 3229 17807 3289 21469
rect 10650 21275 10710 38950
rect 3455 21215 10710 21275
rect 3455 20027 3515 21215
rect 4014 21125 4107 21130
rect 4010 21042 4019 21125
rect 4102 21042 4111 21125
rect 4014 20312 4107 21042
rect 9159 21003 9252 21009
rect 9252 20910 9323 21003
rect 9416 20910 9425 21003
rect 9159 20904 9252 20910
rect 10850 20839 10910 42350
rect 7505 20779 10910 20839
rect 7505 20474 7565 20779
rect 11050 20625 11110 42570
rect 8681 20565 11110 20625
rect 11210 32690 11270 42790
rect 11375 42664 11435 42802
rect 11375 42595 11435 42604
rect 11520 38278 11580 38280
rect 11513 38222 11522 38278
rect 11578 38222 11587 38278
rect 11520 37333 11580 38222
rect 12417 37503 12477 37512
rect 12072 37441 12078 37493
rect 12130 37441 12136 37493
rect 11520 37267 11580 37273
rect 11367 37039 11373 37101
rect 11435 37039 11441 37101
rect 11373 36652 11435 37039
rect 12088 36983 12120 37441
rect 12417 37434 12477 37443
rect 12431 37332 12463 37434
rect 12415 37280 12421 37332
rect 12473 37280 12479 37332
rect 12078 36977 12130 36983
rect 12068 36925 12078 36974
rect 12130 36925 12149 36974
rect 11364 36590 11373 36652
rect 11435 36590 11444 36652
rect 8681 20475 8741 20565
rect 8675 20415 8681 20475
rect 8741 20415 8747 20475
rect 11210 20467 11270 32630
rect 11752 32507 11808 32514
rect 11371 32447 11377 32507
rect 11437 32505 11810 32507
rect 11437 32449 11752 32505
rect 11808 32449 11810 32505
rect 11437 32447 11810 32449
rect 11752 32440 11808 32447
rect 12068 32250 12149 36925
rect 11445 32190 11505 32199
rect 11445 32121 11505 32130
rect 12067 32167 12149 32250
rect 11451 31976 11499 32121
rect 11449 31970 11501 31976
rect 12067 31947 12148 32167
rect 11449 31912 11501 31918
rect 11813 31866 12148 31947
rect 11813 31599 11894 31866
rect 11813 31547 11837 31599
rect 11889 31547 11895 31599
rect 11348 31201 11412 31207
rect 11348 31013 11412 31137
rect 11813 31083 11894 31547
rect 12270 31462 12279 31522
rect 12339 31462 12348 31522
rect 12293 31430 12325 31462
rect 12277 31378 12283 31430
rect 12335 31378 12341 31430
rect 11813 31031 11837 31083
rect 11889 31031 11894 31083
rect 11339 30949 11348 31013
rect 11412 30949 11421 31013
rect 11591 26534 11647 26541
rect 11380 26474 11386 26534
rect 11446 26532 11649 26534
rect 11446 26476 11591 26532
rect 11647 26476 11649 26532
rect 11446 26474 11649 26476
rect 11591 26467 11647 26474
rect 11813 25633 11894 31031
rect 11798 25581 11804 25633
rect 11856 25581 11894 25633
rect 11813 25123 11894 25581
rect 12252 25391 12258 25443
rect 12310 25433 12316 25443
rect 12365 25433 12374 25447
rect 12310 25401 12374 25433
rect 12310 25391 12316 25401
rect 12365 25387 12374 25401
rect 12434 25387 12443 25447
rect 11804 25117 11894 25123
rect 11856 25065 11894 25117
rect 11804 25059 11894 25065
rect 7505 20408 7565 20414
rect 9612 20407 9618 20467
rect 9678 20407 11270 20467
rect 4014 20260 4026 20312
rect 4078 20260 4107 20312
rect 4014 20244 4107 20260
rect 4471 20305 4546 20319
rect 6564 20307 6616 20313
rect 4471 20257 6564 20305
rect 3449 19967 3455 20027
rect 3515 19967 3521 20027
rect 4036 19802 4068 20244
rect 4026 19796 4078 19802
rect 4026 19738 4078 19744
rect 4303 19386 4309 19438
rect 4361 19429 4367 19438
rect 4471 19429 4546 20257
rect 6564 20249 6616 20255
rect 11813 20308 11894 25059
rect 11207 20209 11267 20211
rect 7169 20114 7175 20183
rect 7244 20114 7250 20183
rect 7175 19986 7244 20114
rect 7702 20076 7708 20128
rect 7760 20076 7766 20128
rect 8172 20120 8178 20189
rect 8247 20120 8253 20189
rect 7717 19980 7751 20076
rect 8178 20021 8247 20120
rect 8653 20067 8659 20119
rect 8711 20067 8717 20119
rect 9170 20117 9176 20186
rect 9245 20117 9251 20186
rect 11200 20153 11209 20209
rect 11265 20153 11274 20209
rect 7175 19908 7244 19917
rect 7704 19971 7764 19980
rect 8668 19988 8702 20067
rect 9176 20036 9245 20117
rect 8178 19943 8247 19952
rect 8655 19979 8715 19988
rect 7704 19902 7764 19911
rect 9176 19958 9245 19967
rect 8655 19910 8715 19919
rect 10954 19604 11014 19610
rect 10630 19544 10639 19604
rect 10699 19544 10954 19604
rect 10954 19538 11014 19544
rect 4361 19395 4546 19429
rect 4361 19386 4367 19395
rect 4025 19020 4108 19024
rect 4020 19015 4113 19020
rect 4020 18932 4025 19015
rect 4108 18932 4113 19015
rect 4020 18098 4113 18932
rect 4020 18046 4056 18098
rect 4108 18046 4114 18098
rect 4020 18042 4113 18046
rect 3223 17747 3229 17807
rect 3289 17747 3295 17807
rect 4066 17588 4098 18042
rect 4056 17582 4108 17588
rect 4056 17524 4108 17530
rect 4330 17161 4336 17213
rect 4388 17204 4394 17213
rect 4471 17204 4546 19395
rect 11207 19301 11267 20153
rect 11813 20151 11899 20308
rect 11818 19871 11899 20151
rect 11818 19790 11953 19871
rect 11207 19235 11267 19241
rect 11872 19461 11953 19790
rect 11872 19409 11896 19461
rect 11948 19409 11954 19461
rect 12338 19456 12347 19516
rect 12407 19456 12416 19516
rect 10916 19001 10925 19061
rect 10985 19060 10994 19061
rect 11185 19060 11244 19066
rect 10985 19001 11185 19060
rect 11185 18995 11244 19001
rect 11872 18945 11953 19409
rect 12361 19304 12393 19456
rect 12345 19252 12351 19304
rect 12403 19252 12409 19304
rect 11872 18893 11896 18945
rect 11948 18893 11953 18945
rect 5210 18751 5262 18757
rect 5534 18748 5543 18756
rect 5262 18703 5543 18748
rect 5210 18693 5262 18699
rect 5534 18696 5543 18703
rect 5603 18696 5612 18756
rect 5185 17912 5237 17918
rect 5499 17908 5508 17916
rect 5237 17864 5508 17908
rect 5185 17854 5237 17860
rect 5499 17856 5508 17864
rect 5568 17856 5577 17916
rect 4388 17170 4546 17204
rect 4388 17161 4394 17170
rect 4040 15820 4046 15872
rect 4098 15820 4104 15872
rect 3016 15527 3022 15587
rect 3082 15527 3088 15587
rect 4056 15382 4088 15820
rect 4035 15356 4128 15382
rect 4035 15304 4046 15356
rect 4098 15304 4128 15356
rect 4035 15195 4128 15304
rect 4471 15349 4546 17170
rect 5203 16990 5255 16996
rect 5531 16986 5540 16995
rect 5255 16943 5540 16986
rect 5203 16932 5255 16938
rect 5531 16935 5540 16943
rect 5600 16935 5609 16995
rect 7523 16356 7583 16365
rect 6759 16342 6819 16351
rect 6759 16273 6819 16282
rect 6936 16281 6942 16333
rect 6994 16324 7000 16333
rect 7121 16324 7130 16337
rect 6994 16290 7130 16324
rect 6994 16281 7000 16290
rect 7121 16277 7130 16290
rect 7190 16277 7199 16337
rect 7523 16287 7583 16296
rect 8057 16347 8109 16353
rect 8309 16351 8369 16360
rect 8109 16304 8309 16338
rect 8057 16289 8109 16295
rect 6759 16122 6818 16273
rect 7523 16094 7582 16287
rect 8309 16282 8369 16291
rect 8922 16343 8982 16352
rect 8922 16274 8982 16283
rect 8922 16113 8981 16274
rect 6759 16057 6818 16063
rect 7517 16035 7523 16094
rect 7582 16035 7588 16094
rect 8916 16054 8922 16113
rect 8981 16054 8987 16113
rect 5049 15515 5055 15575
rect 5115 15515 5121 15575
rect 4596 15349 4602 15358
rect 4471 15315 4602 15349
rect 4471 15290 4546 15315
rect 4596 15306 4602 15315
rect 4654 15306 4660 15358
rect 4035 15112 4040 15195
rect 4123 15112 4128 15195
rect 4035 15107 4128 15112
rect 4040 15103 4123 15107
rect 5055 14922 5115 15515
rect 6601 15498 6607 15558
rect 6667 15498 6673 15558
rect 2794 14862 5115 14922
rect 6013 15349 6106 15355
rect 6013 14878 6106 15256
rect 6009 14795 6018 14878
rect 6101 14795 6110 14878
rect 6013 14790 6106 14795
rect 6607 14675 6667 15498
rect 8054 15488 8060 15548
rect 8120 15488 8126 15548
rect 2582 14615 6667 14675
rect 8060 14350 8120 15488
rect 9134 15372 9143 15434
rect 9205 15372 9214 15434
rect 8676 15318 8738 15324
rect 9143 15318 9205 15372
rect 8738 15256 9205 15318
rect 8676 15250 8738 15256
rect 11872 14361 11953 18893
rect 2323 14290 8120 14350
rect 11172 14305 11232 14307
rect 11165 14249 11174 14305
rect 11230 14249 11239 14305
rect 7625 13941 7718 13947
rect 5020 13501 5029 13561
rect 5089 13560 5098 13561
rect 5530 13560 5588 13566
rect 5089 13502 5530 13560
rect 5089 13501 5098 13502
rect 5530 13496 5588 13502
rect 7625 8258 7718 13848
rect 10532 13654 10593 13663
rect 10824 13654 10885 13660
rect 10593 13593 10824 13654
rect 10532 13584 10593 13593
rect 10824 13587 10885 13593
rect 11172 13349 11232 14249
rect 11870 14247 11953 14361
rect 11870 13883 11951 14247
rect 11172 13283 11232 13289
rect 11765 13802 11951 13883
rect 11765 13508 11846 13802
rect 11765 13456 11796 13508
rect 11848 13456 11854 13508
rect 12359 13466 12368 13526
rect 12428 13466 12437 13526
rect 10835 13058 10844 13118
rect 10904 13117 10913 13118
rect 11156 13117 11214 13123
rect 10904 13059 11156 13117
rect 10904 13058 10913 13059
rect 11156 13053 11214 13059
rect 11765 12998 11846 13456
rect 12238 13345 12290 13351
rect 12382 13335 12414 13466
rect 12290 13303 12414 13335
rect 12238 13287 12290 13293
rect 11765 12992 11848 12998
rect 11765 12940 11796 12992
rect 11765 12934 11848 12940
rect 11185 8377 11241 8384
rect 11183 8375 11243 8377
rect 11183 8319 11185 8375
rect 11241 8319 11243 8375
rect 7621 8175 7630 8258
rect 7713 8175 7722 8258
rect 7625 8170 7718 8175
rect 10942 7759 11007 7765
rect 10675 7694 10684 7759
rect 10749 7694 10942 7759
rect 10942 7688 11007 7694
rect 11183 7440 11243 8319
rect 11765 7609 11846 12934
rect 11764 7557 11770 7609
rect 11822 7557 11846 7609
rect 11183 7374 11243 7380
rect 11182 7215 11243 7221
rect 10864 7154 10873 7215
rect 10934 7154 11182 7215
rect 11182 7148 11243 7154
rect 11765 7093 11846 7557
rect 12355 7453 12364 7513
rect 12424 7453 12433 7513
rect 12238 7398 12290 7404
rect 12378 7388 12410 7453
rect 12290 7356 12410 7388
rect 12238 7340 12290 7346
rect 11765 7041 11770 7093
rect 11822 7041 11846 7093
rect 11765 2685 11846 7041
rect 11765 2604 12036 2685
rect 11375 1438 11435 1440
rect 10911 1356 10920 1416
rect 10980 1415 10989 1416
rect 11177 1415 11236 1421
rect 10980 1356 11177 1415
rect 11368 1382 11377 1438
rect 11433 1382 11442 1438
rect 11177 1350 11236 1356
rect 11375 1111 11435 1382
rect 11955 1266 12036 2604
rect 12396 1386 12462 1391
rect 12392 1330 12401 1386
rect 12457 1330 12466 1386
rect 11955 1214 11976 1266
rect 12028 1214 12036 1266
rect 11955 1194 12036 1214
rect 11375 1045 11435 1051
rect 11367 860 11427 866
rect 11137 800 11146 860
rect 11206 800 11367 860
rect 11367 794 11427 800
rect 11986 787 12018 1194
rect 12396 1150 12462 1330
rect 12396 1078 12462 1084
rect 30515 830 30685 834
rect 12486 825 30690 830
rect 12486 787 30515 825
rect 11965 750 30515 787
rect 11965 698 11976 750
rect 12028 698 30515 750
rect 11965 694 30515 698
rect 11976 692 12028 694
rect 12486 655 30515 694
rect 30685 655 30690 825
rect 12486 650 30690 655
rect 30515 646 30685 650
<< via2 >>
rect 9352 44712 9408 44768
rect 6632 44092 6688 44148
rect 8294 44080 8354 44140
rect 3152 43672 3208 43728
rect 9752 44532 9808 44588
rect 11840 44552 11896 44608
rect 12576 44572 12632 44628
rect 9350 43590 9410 43650
rect 9130 42570 9190 42630
rect 9290 42350 9350 42410
rect 9370 38950 9430 39010
rect 950 37610 1010 37670
rect 770 34210 830 34270
rect 1130 36230 1190 36290
rect 9430 34870 9490 34930
rect 9352 33932 9408 33988
rect 5472 33132 5528 33188
rect 9555 32864 9625 32934
rect 9634 32437 9690 32493
rect 13312 44552 13368 44608
rect 14048 44572 14104 44628
rect 14784 44572 14840 44628
rect 9920 32435 9980 32495
rect 9269 26688 9334 26753
rect 9555 25379 9615 25439
rect 8167 24241 8250 24324
rect 7166 23909 7249 23992
rect 1659 20391 1736 20468
rect 1673 18184 1733 18244
rect 1692 15956 1752 16016
rect 15520 44552 15576 44608
rect 16256 44552 16312 44608
rect 24352 44601 24408 44657
rect 16992 44512 17048 44568
rect 4019 21042 4102 21125
rect 9323 20910 9416 21003
rect 11375 42604 11435 42664
rect 11522 38222 11578 38278
rect 12417 37443 12477 37503
rect 11373 36590 11435 36652
rect 11752 32449 11808 32505
rect 11445 32130 11505 32190
rect 12279 31462 12339 31522
rect 11348 30949 11412 31013
rect 11591 26476 11647 26532
rect 12374 25387 12434 25447
rect 7175 19917 7244 19986
rect 11209 20153 11265 20209
rect 7704 19911 7764 19971
rect 8178 19952 8247 20021
rect 8655 19919 8715 19979
rect 9176 19967 9245 20036
rect 10639 19544 10699 19604
rect 4025 18932 4108 19015
rect 12347 19456 12407 19516
rect 10925 19001 10985 19061
rect 5543 18696 5603 18756
rect 5508 17856 5568 17916
rect 5540 16935 5600 16995
rect 6759 16282 6819 16342
rect 7130 16277 7190 16337
rect 7523 16296 7583 16356
rect 8309 16291 8369 16351
rect 8922 16283 8982 16343
rect 4040 15112 4123 15195
rect 6018 14795 6101 14878
rect 9143 15372 9205 15434
rect 11174 14249 11230 14305
rect 5029 13501 5089 13561
rect 10532 13593 10593 13654
rect 12368 13466 12428 13526
rect 10844 13058 10904 13118
rect 11185 8319 11241 8375
rect 7630 8175 7713 8258
rect 10684 7694 10749 7759
rect 10873 7154 10934 7215
rect 12364 7453 12424 7513
rect 10920 1356 10980 1416
rect 11377 1382 11433 1438
rect 12401 1330 12457 1386
rect 11146 800 11206 860
rect 30515 655 30685 825
<< metal3 >>
rect 9347 44770 9413 44773
rect 10364 44772 10428 44778
rect 9347 44768 10364 44770
rect 8156 44752 8220 44758
rect 390 44690 8156 44750
rect 390 33190 450 44690
rect 9347 44712 9352 44768
rect 9408 44712 10364 44768
rect 9347 44710 10364 44712
rect 9347 44707 9413 44710
rect 11094 44728 11100 44792
rect 11164 44728 11170 44792
rect 11830 44728 11836 44792
rect 11900 44728 11906 44792
rect 12566 44748 12572 44812
rect 12636 44748 12642 44812
rect 13302 44748 13308 44812
rect 13372 44748 13378 44812
rect 14038 44748 14044 44812
rect 14108 44748 14114 44812
rect 10364 44702 10428 44708
rect 8156 44682 8220 44688
rect 988 44592 1052 44598
rect 610 44530 988 44590
rect 610 43050 670 44530
rect 988 44522 1052 44528
rect 9747 44590 9813 44593
rect 11102 44590 11162 44728
rect 11838 44613 11898 44728
rect 12574 44633 12634 44748
rect 12571 44628 12637 44633
rect 9747 44588 11162 44590
rect 9747 44532 9752 44588
rect 9808 44532 11162 44588
rect 11835 44608 11901 44613
rect 11835 44552 11840 44608
rect 11896 44552 11901 44608
rect 12571 44572 12576 44628
rect 12632 44572 12637 44628
rect 13310 44613 13370 44748
rect 14046 44633 14106 44748
rect 14774 44728 14780 44792
rect 14844 44728 14850 44792
rect 15510 44748 15516 44812
rect 15580 44748 15586 44812
rect 14782 44633 14842 44728
rect 14043 44628 14109 44633
rect 12571 44567 12637 44572
rect 13307 44608 13373 44613
rect 11835 44547 11901 44552
rect 13307 44552 13312 44608
rect 13368 44552 13373 44608
rect 14043 44572 14048 44628
rect 14104 44572 14109 44628
rect 14043 44567 14109 44572
rect 14779 44628 14845 44633
rect 14779 44572 14784 44628
rect 14840 44572 14845 44628
rect 15518 44613 15578 44748
rect 16246 44708 16252 44772
rect 16316 44708 16322 44772
rect 16982 44728 16988 44792
rect 17052 44728 17058 44792
rect 24342 44749 24348 44813
rect 24412 44749 24418 44813
rect 16254 44613 16314 44708
rect 14779 44567 14845 44572
rect 15515 44608 15581 44613
rect 13307 44547 13373 44552
rect 15515 44552 15520 44608
rect 15576 44552 15581 44608
rect 15515 44547 15581 44552
rect 16251 44608 16317 44613
rect 16251 44552 16256 44608
rect 16312 44552 16317 44608
rect 16990 44573 17050 44728
rect 24350 44662 24410 44749
rect 24347 44657 24413 44662
rect 24347 44601 24352 44657
rect 24408 44601 24413 44657
rect 24347 44596 24413 44601
rect 16251 44547 16317 44552
rect 16987 44568 17053 44573
rect 9747 44530 11162 44532
rect 9747 44527 9813 44530
rect 16987 44512 16992 44568
rect 17048 44512 17053 44568
rect 16987 44507 17053 44512
rect 30971 44404 31035 44410
rect 8294 44342 30971 44402
rect 6627 44150 6693 44153
rect 8068 44152 8132 44158
rect 6627 44148 8068 44150
rect 6627 44092 6632 44148
rect 6688 44092 8068 44148
rect 6627 44090 8068 44092
rect 6627 44087 6693 44090
rect 8294 44145 8354 44342
rect 30971 44334 31035 44340
rect 8068 44082 8132 44088
rect 8289 44140 8359 44145
rect 8289 44080 8294 44140
rect 8354 44080 8359 44140
rect 22401 44086 22465 44092
rect 8289 44075 8359 44080
rect 20899 44024 22401 44084
rect 3147 43730 3213 43733
rect 3147 43728 3650 43730
rect 3147 43672 3152 43728
rect 3208 43672 3650 43728
rect 3147 43670 3650 43672
rect 3147 43667 3213 43670
rect 3590 42630 3650 43670
rect 9345 43650 9415 43655
rect 9345 43590 9350 43650
rect 9410 43590 9415 43650
rect 9345 43585 9415 43590
rect 9350 43418 9410 43585
rect 9348 43412 9412 43418
rect 9348 43342 9412 43348
rect 11564 43223 11570 43287
rect 11634 43285 11640 43287
rect 20899 43285 20959 44024
rect 22401 44016 22465 44022
rect 22413 43926 22477 43932
rect 11634 43225 20959 43285
rect 21071 43864 22413 43924
rect 11634 43223 11640 43225
rect 11732 43010 11738 43074
rect 11802 43072 11808 43074
rect 21071 43072 21131 43864
rect 22413 43856 22477 43862
rect 21278 43755 21342 43761
rect 22405 43755 22469 43761
rect 21342 43693 22405 43753
rect 21278 43685 21342 43691
rect 22405 43685 22469 43691
rect 22392 43545 22456 43551
rect 21438 43481 21444 43545
rect 21508 43543 21514 43545
rect 21508 43483 22392 43543
rect 21508 43481 21514 43483
rect 22392 43475 22456 43481
rect 22387 43291 22451 43297
rect 21615 43227 21621 43291
rect 21685 43289 21691 43291
rect 21685 43229 22387 43289
rect 21685 43227 21691 43229
rect 22387 43221 22451 43227
rect 11802 43012 21131 43072
rect 22393 43061 22457 43067
rect 11802 43010 11808 43012
rect 21796 42997 21802 43061
rect 21866 43059 21872 43061
rect 21866 42999 22393 43059
rect 21866 42997 21872 42999
rect 22393 42991 22457 42997
rect 10383 42901 10507 42913
rect 22404 42901 22499 42906
rect 10383 42900 22500 42901
rect 10383 42805 22404 42900
rect 22499 42805 22500 42900
rect 10383 42804 22500 42805
rect 10383 42716 10511 42804
rect 22404 42799 22499 42804
rect 9125 42630 9195 42635
rect 3590 42570 9130 42630
rect 9190 42570 9195 42630
rect 9125 42565 9195 42570
rect 9285 42410 9355 42415
rect 9150 42350 9290 42410
rect 9350 42350 9355 42410
rect 9285 42345 9355 42350
rect 1222 41730 1228 41732
rect 1090 41670 1228 41730
rect 1222 41668 1228 41670
rect 1292 41668 1298 41732
rect 982 39948 988 40012
rect 1052 39948 1058 40012
rect 990 39650 1050 39948
rect 9365 39010 9435 39015
rect 9270 38950 9370 39010
rect 9430 38950 9435 39010
rect 9365 38945 9435 38950
rect 945 37670 1015 37675
rect 770 37610 950 37670
rect 1010 37610 1015 37670
rect 945 37605 1015 37610
rect 10383 37008 10507 42716
rect 11370 42664 11440 42669
rect 11370 42604 11375 42664
rect 11435 42604 11440 42664
rect 11370 42599 11440 42604
rect 11375 42448 11435 42599
rect 11373 42442 11437 42448
rect 11373 42372 11437 42378
rect 9631 36888 10507 37008
rect 10383 36886 10507 36888
rect 10741 39353 13307 39446
rect 1125 36290 1195 36295
rect 870 36230 1130 36290
rect 1190 36230 1195 36290
rect 1125 36225 1195 36230
rect 9425 34930 9495 34935
rect 9310 34870 9430 34930
rect 9490 34870 9495 34930
rect 9425 34865 9495 34870
rect 9342 34628 9348 34692
rect 9412 34628 9418 34692
rect 765 34270 835 34275
rect 765 34210 770 34270
rect 830 34210 990 34270
rect 765 34205 835 34210
rect 9350 33993 9410 34628
rect 9347 33988 9413 33993
rect 9347 33932 9352 33988
rect 9408 33932 9413 33988
rect 9347 33927 9413 33932
rect 5467 33190 5533 33193
rect 390 33188 5533 33190
rect 390 33132 5472 33188
rect 5528 33132 5533 33188
rect 390 33130 5533 33132
rect 5467 33127 5533 33130
rect 9550 32934 9630 32939
rect 9296 32864 9302 32934
rect 9372 32864 9555 32934
rect 9625 32864 9630 32934
rect 9550 32859 9630 32864
rect 9629 32495 9695 32498
rect 9915 32495 9985 32500
rect 9629 32493 9920 32495
rect 9629 32437 9634 32493
rect 9690 32437 9920 32493
rect 9629 32435 9920 32437
rect 9980 32435 9985 32495
rect 9629 32432 9695 32435
rect 9915 32430 9985 32435
rect 10265 32192 10329 32198
rect 9564 32128 9570 32192
rect 9634 32190 9640 32192
rect 9634 32130 10265 32190
rect 9634 32128 9640 32130
rect 10265 32122 10329 32128
rect 9264 26753 9339 26758
rect 8988 26688 8994 26753
rect 9059 26688 9269 26753
rect 9334 26688 9339 26753
rect 9264 26683 9339 26688
rect 9553 25666 9617 25672
rect 9553 25596 9617 25602
rect 9555 25444 9615 25596
rect 9550 25439 9620 25444
rect 9550 25379 9555 25439
rect 9615 25379 9620 25439
rect 9550 25374 9620 25379
rect 10741 24329 10834 39353
rect 11517 38280 11583 38283
rect 12412 38282 12476 38288
rect 11517 38278 12412 38280
rect 11517 38222 11522 38278
rect 11578 38222 12412 38278
rect 11517 38220 12412 38222
rect 11517 38217 11583 38220
rect 12412 38212 12476 38218
rect 12415 37508 12880 37540
rect 12412 37503 12880 37508
rect 12412 37443 12417 37503
rect 12477 37443 12880 37503
rect 12412 37440 12880 37443
rect 12412 37438 12482 37440
rect 10969 36589 10975 36653
rect 11039 36652 11045 36653
rect 11368 36652 11440 36657
rect 11039 36590 11373 36652
rect 11435 36590 11440 36652
rect 11039 36589 11045 36590
rect 11368 36585 11440 36590
rect 8162 24324 10834 24329
rect 8162 24241 8167 24324
rect 8250 24241 10834 24324
rect 8162 24236 10834 24241
rect 10975 33634 13296 33727
rect 10975 23997 11068 33634
rect 11747 32507 11813 32510
rect 12249 32509 12313 32515
rect 11747 32505 12249 32507
rect 11747 32449 11752 32505
rect 11808 32449 12249 32505
rect 11747 32447 12249 32449
rect 11747 32444 11813 32447
rect 12249 32439 12313 32445
rect 11199 32128 11205 32192
rect 11269 32190 11275 32192
rect 11440 32190 11510 32195
rect 11269 32130 11445 32190
rect 11505 32130 11510 32190
rect 11269 32128 11275 32130
rect 11440 32125 11510 32130
rect 12274 31522 12344 31527
rect 12548 31522 12780 31540
rect 12274 31462 12279 31522
rect 12339 31462 12780 31522
rect 12274 31457 12344 31462
rect 12548 31440 12780 31462
rect 11343 31013 11417 31018
rect 11182 30949 11188 31013
rect 11252 30949 11348 31013
rect 11412 30949 11417 31013
rect 11343 30944 11417 30949
rect 7161 23992 11068 23997
rect 7161 23909 7166 23992
rect 7249 23909 11068 23992
rect 7161 23904 11068 23909
rect 11193 27271 13318 27364
rect 11193 23707 11286 27271
rect 11586 26534 11652 26537
rect 12085 26536 12149 26542
rect 11586 26532 12085 26534
rect 11586 26476 11591 26532
rect 11647 26476 12085 26532
rect 11586 26474 12085 26476
rect 11586 26471 11652 26474
rect 12085 26466 12149 26472
rect 12374 25540 12434 25548
rect 12374 25452 12840 25540
rect 12369 25447 12840 25452
rect 12369 25387 12374 25447
rect 12434 25440 12840 25447
rect 12434 25387 12439 25440
rect 12369 25382 12439 25387
rect 4014 23614 11286 23707
rect 4014 21125 4107 23614
rect 4014 21042 4019 21125
rect 4102 21042 4107 21125
rect 4014 21037 4107 21042
rect 4567 21161 13263 21254
rect 1654 20468 1741 20473
rect 1275 20391 1281 20468
rect 1358 20391 1659 20468
rect 1736 20391 1741 20468
rect 1654 20386 1741 20391
rect 4567 19020 4660 21161
rect 9318 21003 9421 21008
rect 9318 20910 9323 21003
rect 9416 20910 9514 21003
rect 9607 20910 9613 21003
rect 9318 20905 9421 20910
rect 11204 20211 11270 20214
rect 11925 20213 11989 20219
rect 11204 20209 11925 20211
rect 11204 20153 11209 20209
rect 11265 20153 11925 20209
rect 11204 20151 11925 20153
rect 11204 20148 11270 20151
rect 11925 20143 11989 20149
rect 9171 20036 9250 20041
rect 8173 20021 8252 20026
rect 7170 19986 7249 19991
rect 7170 19917 7175 19986
rect 7244 19917 7249 19986
rect 7170 19912 7249 19917
rect 7699 19971 7769 19976
rect 7852 19971 7858 19973
rect 7175 19399 7244 19912
rect 7699 19911 7704 19971
rect 7764 19911 7858 19971
rect 7699 19906 7769 19911
rect 7852 19909 7858 19911
rect 7922 19909 7928 19973
rect 8173 19952 8178 20021
rect 8247 19952 8252 20021
rect 8173 19947 8252 19952
rect 8650 19979 8720 19984
rect 8831 19979 8837 19981
rect 8178 19417 8247 19947
rect 8650 19919 8655 19979
rect 8715 19919 8837 19979
rect 8650 19914 8720 19919
rect 8831 19917 8837 19919
rect 8901 19917 8907 19981
rect 9171 19967 9176 20036
rect 9245 19967 9250 20036
rect 9171 19962 9250 19967
rect 9176 19402 9245 19962
rect 10634 19604 10704 19609
rect 10373 19544 10639 19604
rect 10699 19544 10704 19604
rect 4020 19015 4660 19020
rect 4020 18932 4025 19015
rect 4108 18932 4660 19015
rect 4020 18927 4660 18932
rect 5538 18756 5608 18761
rect 5538 18696 5543 18756
rect 5603 18696 6717 18756
rect 10373 18728 10433 19544
rect 10634 19539 10704 19544
rect 12548 19521 12840 19540
rect 12342 19516 12840 19521
rect 12342 19456 12347 19516
rect 12407 19456 12840 19516
rect 12342 19451 12840 19456
rect 12548 19440 12840 19451
rect 10632 18999 10638 19063
rect 10702 19061 10708 19063
rect 10920 19061 10990 19066
rect 10702 19001 10925 19061
rect 10985 19001 10990 19061
rect 10702 18999 10708 19001
rect 10920 18996 10990 19001
rect 10371 18722 10435 18728
rect 5538 18691 5608 18696
rect 10371 18652 10435 18658
rect 1287 18182 1293 18246
rect 1357 18244 1363 18246
rect 1668 18244 1738 18249
rect 1357 18184 1673 18244
rect 1733 18184 1738 18244
rect 1357 18182 1363 18184
rect 1668 18179 1738 18184
rect 5503 17916 5573 17921
rect 5503 17856 5508 17916
rect 5568 17856 6735 17916
rect 5503 17851 5573 17856
rect 5535 16995 5605 17000
rect 5535 16935 5540 16995
rect 5600 16935 6837 16995
rect 5535 16930 5605 16935
rect 6759 16347 6819 16906
rect 7523 16361 7583 16985
rect 7518 16356 7588 16361
rect 6754 16342 6824 16347
rect 6754 16282 6759 16342
rect 6819 16282 6824 16342
rect 6754 16277 6824 16282
rect 7125 16337 7195 16342
rect 7125 16277 7130 16337
rect 7190 16277 7195 16337
rect 7518 16296 7523 16356
rect 7583 16296 7588 16356
rect 7518 16291 7588 16296
rect 8304 16351 8374 16356
rect 8304 16291 8309 16351
rect 8369 16291 8374 16351
rect 8922 16348 8982 17008
rect 8304 16286 8374 16291
rect 8917 16343 8987 16348
rect 7125 16272 7195 16277
rect 7130 16196 7190 16272
rect 8309 16203 8369 16286
rect 8917 16283 8922 16343
rect 8982 16283 8987 16343
rect 8917 16278 8987 16283
rect 8307 16197 8371 16203
rect 7128 16190 7192 16196
rect 8307 16127 8371 16133
rect 7128 16120 7192 16126
rect 1335 15954 1341 16018
rect 1405 16016 1411 16018
rect 1687 16016 1757 16021
rect 1405 15956 1692 16016
rect 1752 15956 1757 16016
rect 1405 15954 1411 15956
rect 1687 15951 1757 15956
rect 9138 15434 9210 15439
rect 9359 15434 9365 15435
rect 9138 15372 9143 15434
rect 9205 15372 9365 15434
rect 9138 15367 9210 15372
rect 9359 15371 9365 15372
rect 9429 15371 9435 15435
rect 4035 15195 13312 15200
rect 4035 15112 4040 15195
rect 4123 15112 13312 15195
rect 4035 15107 13312 15112
rect 6013 14878 6106 14883
rect 6013 14795 6018 14878
rect 6101 14795 6106 14878
rect 865 13499 871 13563
rect 935 13561 941 13563
rect 5024 13561 5094 13566
rect 935 13501 5029 13561
rect 5089 13501 5094 13561
rect 935 13499 941 13501
rect 5024 13496 5094 13501
rect 6013 8748 6106 14795
rect 9121 14398 9419 14403
rect 9120 14397 10389 14398
rect 9120 14099 9121 14397
rect 9419 14099 10389 14397
rect 9120 14098 10389 14099
rect 10689 14098 10695 14398
rect 11169 14307 11235 14310
rect 11738 14309 11802 14315
rect 11169 14305 11738 14307
rect 11169 14249 11174 14305
rect 11230 14249 11738 14305
rect 11169 14247 11738 14249
rect 11169 14244 11235 14247
rect 11738 14239 11802 14245
rect 9121 14093 9419 14098
rect 10531 13903 10595 13909
rect 10531 13833 10595 13839
rect 10532 13659 10593 13833
rect 10527 13654 10598 13659
rect 10527 13593 10532 13654
rect 10593 13593 10598 13654
rect 10527 13588 10598 13593
rect 12537 13539 12820 13540
rect 12356 13526 12820 13539
rect 12356 13466 12368 13526
rect 12428 13466 12820 13526
rect 12356 13454 12820 13466
rect 12537 13440 12820 13454
rect 10474 13056 10480 13120
rect 10544 13118 10550 13120
rect 10839 13118 10909 13123
rect 10544 13058 10844 13118
rect 10904 13058 10909 13118
rect 10544 13056 10550 13058
rect 10839 13053 10909 13058
rect 6013 8655 13346 8748
rect 11180 8377 11246 8380
rect 11570 8379 11634 8385
rect 11180 8375 11570 8377
rect 11180 8319 11185 8375
rect 11241 8319 11570 8375
rect 11180 8317 11570 8319
rect 11180 8314 11246 8317
rect 11570 8309 11634 8315
rect 7625 8258 7718 8263
rect 7625 8175 7630 8258
rect 7713 8175 7718 8258
rect 7625 3808 7718 8175
rect 10679 7759 10754 7764
rect 9599 7694 9605 7759
rect 9670 7694 10684 7759
rect 10749 7694 10754 7759
rect 10679 7689 10754 7694
rect 12349 7513 12820 7540
rect 12349 7453 12364 7513
rect 12424 7453 12820 7513
rect 12349 7440 12820 7453
rect 10502 7153 10508 7217
rect 10572 7215 10578 7217
rect 10868 7215 10939 7220
rect 10572 7154 10873 7215
rect 10934 7154 10939 7215
rect 10572 7153 10578 7154
rect 10868 7149 10939 7154
rect 7625 3715 13274 3808
rect 11367 1570 11373 1634
rect 11437 1570 11443 1634
rect 11375 1443 11435 1570
rect 11372 1438 11438 1443
rect 12379 1440 12800 1540
rect 9329 1418 9393 1424
rect 10915 1416 10985 1421
rect 9393 1356 10920 1416
rect 10980 1356 10985 1416
rect 11372 1382 11377 1438
rect 11433 1382 11438 1438
rect 11372 1377 11438 1382
rect 12396 1386 12462 1440
rect 9329 1348 9393 1354
rect 10915 1351 10985 1356
rect 12396 1330 12401 1386
rect 12457 1330 12462 1386
rect 12396 1325 12462 1330
rect 10923 798 10929 862
rect 10993 860 10999 862
rect 11141 860 11211 865
rect 10993 800 11146 860
rect 11206 800 11211 860
rect 10993 798 10999 800
rect 11141 795 11211 800
rect 30510 829 31462 830
rect 30510 825 31283 829
rect 30510 655 30515 825
rect 30685 655 31283 825
rect 30510 651 31283 655
rect 31461 651 31467 829
rect 30510 650 31462 651
<< via3 >>
rect 8156 44688 8220 44752
rect 10364 44708 10428 44772
rect 11100 44728 11164 44792
rect 11836 44728 11900 44792
rect 12572 44748 12636 44812
rect 13308 44748 13372 44812
rect 14044 44748 14108 44812
rect 988 44528 1052 44592
rect 14780 44728 14844 44792
rect 15516 44748 15580 44812
rect 16252 44708 16316 44772
rect 16988 44728 17052 44792
rect 24348 44749 24412 44813
rect 8068 44088 8132 44152
rect 30971 44340 31035 44404
rect 9348 43348 9412 43412
rect 11570 43223 11634 43287
rect 22401 44022 22465 44086
rect 11738 43010 11802 43074
rect 22413 43862 22477 43926
rect 21278 43691 21342 43755
rect 22405 43691 22469 43755
rect 21444 43481 21508 43545
rect 22392 43481 22456 43545
rect 21621 43227 21685 43291
rect 22387 43227 22451 43291
rect 21802 42997 21866 43061
rect 22393 42997 22457 43061
rect 22404 42805 22499 42900
rect 1228 41668 1292 41732
rect 988 39948 1052 40012
rect 11373 42378 11437 42442
rect 9348 34628 9412 34692
rect 9302 32864 9372 32934
rect 9570 32128 9634 32192
rect 10265 32128 10329 32192
rect 8994 26688 9059 26753
rect 9553 25602 9617 25666
rect 12412 38218 12476 38282
rect 10975 36589 11039 36653
rect 12249 32445 12313 32509
rect 11205 32128 11269 32192
rect 11188 30949 11252 31013
rect 12085 26472 12149 26536
rect 1281 20391 1358 20468
rect 9514 20910 9607 21003
rect 11925 20149 11989 20213
rect 7858 19909 7922 19973
rect 8837 19917 8901 19981
rect 10638 18999 10702 19063
rect 10371 18658 10435 18722
rect 1293 18182 1357 18246
rect 7128 16126 7192 16190
rect 8307 16133 8371 16197
rect 1341 15954 1405 16018
rect 9365 15371 9429 15435
rect 871 13499 935 13563
rect 9121 14099 9419 14397
rect 10389 14098 10689 14398
rect 11738 14245 11802 14309
rect 10531 13839 10595 13903
rect 10480 13056 10544 13120
rect 11570 8315 11634 8379
rect 9605 7694 9670 7759
rect 10508 7153 10572 7217
rect 11373 1570 11437 1634
rect 9329 1354 9393 1418
rect 10929 798 10993 862
rect 31283 651 31461 829
<< metal4 >>
rect 798 44773 858 45152
rect 1534 44773 1594 45152
rect 2270 44773 2330 45152
rect 3006 44773 3066 45152
rect 3742 44773 3802 45152
rect 4478 44773 4538 45152
rect 5214 44773 5274 45152
rect 5950 44773 6010 45152
rect 798 44713 6010 44773
rect 200 44050 500 44152
rect 798 44050 858 44713
rect 987 44592 1053 44593
rect 987 44528 988 44592
rect 1052 44590 1053 44592
rect 6686 44590 6746 45152
rect 1052 44530 6746 44590
rect 1052 44528 1053 44530
rect 987 44527 1053 44528
rect 7422 44430 7482 45152
rect 8158 44753 8218 45152
rect 8155 44752 8221 44753
rect 8155 44688 8156 44752
rect 8220 44688 8221 44752
rect 8155 44687 8221 44688
rect 200 43990 858 44050
rect 990 44370 7482 44430
rect 200 34800 500 43990
rect 990 40013 1050 44370
rect 8067 44152 8133 44153
rect 8067 44088 8068 44152
rect 8132 44150 8133 44152
rect 8894 44150 8954 45152
rect 8132 44090 8954 44150
rect 8132 44088 8133 44090
rect 8067 44087 8133 44088
rect 9630 43890 9690 45152
rect 10366 44773 10426 45152
rect 11102 44793 11162 45152
rect 11838 44793 11898 45152
rect 12574 44813 12634 45152
rect 13310 44813 13370 45152
rect 14046 44813 14106 45152
rect 12571 44812 12637 44813
rect 11099 44792 11165 44793
rect 10363 44772 10429 44773
rect 10363 44708 10364 44772
rect 10428 44708 10429 44772
rect 11099 44728 11100 44792
rect 11164 44728 11165 44792
rect 11099 44727 11165 44728
rect 11835 44792 11901 44793
rect 11835 44728 11836 44792
rect 11900 44728 11901 44792
rect 12571 44748 12572 44812
rect 12636 44748 12637 44812
rect 12571 44747 12637 44748
rect 13307 44812 13373 44813
rect 13307 44748 13308 44812
rect 13372 44748 13373 44812
rect 13307 44747 13373 44748
rect 14043 44812 14109 44813
rect 14043 44748 14044 44812
rect 14108 44748 14109 44812
rect 14782 44793 14842 45152
rect 15518 44813 15578 45152
rect 15515 44812 15581 44813
rect 14043 44747 14109 44748
rect 14779 44792 14845 44793
rect 11835 44727 11901 44728
rect 14779 44728 14780 44792
rect 14844 44728 14845 44792
rect 15515 44748 15516 44812
rect 15580 44748 15581 44812
rect 16254 44773 16314 45152
rect 16990 44793 17050 45152
rect 16987 44792 17053 44793
rect 15515 44747 15581 44748
rect 16251 44772 16317 44773
rect 14779 44727 14845 44728
rect 10363 44707 10429 44708
rect 16251 44708 16252 44772
rect 16316 44708 16317 44772
rect 16987 44728 16988 44792
rect 17052 44728 17053 44792
rect 16987 44727 17053 44728
rect 16251 44707 16317 44708
rect 17726 44200 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44814 24410 45152
rect 24347 44813 24413 44814
rect 24347 44749 24348 44813
rect 24412 44749 24413 44813
rect 24347 44748 24413 44749
rect 1230 43830 9690 43890
rect 9800 43853 22293 44200
rect 22400 44086 22466 44087
rect 22400 44022 22401 44086
rect 22465 44084 22466 44086
rect 25086 44084 25146 45152
rect 22465 44024 25146 44084
rect 22465 44022 22466 44024
rect 22400 44021 22466 44022
rect 22412 43926 22478 43927
rect 22412 43862 22413 43926
rect 22477 43924 22478 43926
rect 25822 43924 25882 45152
rect 22477 43864 25882 43924
rect 22477 43862 22478 43864
rect 22412 43861 22478 43862
rect 1230 41733 1290 43830
rect 9800 43600 10122 43853
rect 21277 43755 21343 43756
rect 21277 43691 21278 43755
rect 21342 43691 21343 43755
rect 21277 43690 21343 43691
rect 9347 43412 9413 43413
rect 9347 43348 9348 43412
rect 9412 43348 9413 43412
rect 9347 43347 9413 43348
rect 1227 41732 1293 41733
rect 1227 41668 1228 41732
rect 1292 41668 1293 41732
rect 1227 41667 1293 41668
rect 987 40012 1053 40013
rect 987 39948 988 40012
rect 1052 39948 1053 40012
rect 987 39947 1053 39948
rect 2400 34800 2700 35100
rect 200 34500 2700 34800
rect 8293 34505 8570 35267
rect 9350 34693 9410 43347
rect 9800 36652 10100 43600
rect 21280 43471 21340 43690
rect 21443 43545 21509 43546
rect 21443 43481 21444 43545
rect 21508 43481 21509 43545
rect 21443 43480 21509 43481
rect 11927 43411 21340 43471
rect 11569 43287 11635 43288
rect 11569 43223 11570 43287
rect 11634 43223 11635 43287
rect 11569 43222 11635 43223
rect 11372 42442 11438 42443
rect 11372 42378 11373 42442
rect 11437 42378 11438 42442
rect 11372 42377 11438 42378
rect 10974 36653 11040 36654
rect 10974 36652 10975 36653
rect 9800 36590 10975 36652
rect 9347 34692 9413 34693
rect 9347 34628 9348 34692
rect 9412 34628 9413 34692
rect 9347 34627 9413 34628
rect 9800 34505 10100 36590
rect 10974 36589 10975 36590
rect 11039 36589 11040 36653
rect 10974 36588 11040 36589
rect 200 26193 500 34500
rect 8293 34187 10100 34505
rect 9142 32934 9442 33827
rect 9142 32864 9302 32934
rect 9372 32864 9442 32934
rect 9142 32190 9442 32864
rect 9569 32192 9635 32193
rect 9569 32190 9570 32192
rect 9142 32130 9570 32190
rect 8993 26753 9060 26754
rect 9142 26753 9442 32130
rect 9569 32128 9570 32130
rect 9634 32128 9635 32192
rect 9569 32127 9635 32128
rect 8993 26688 8994 26753
rect 9059 26688 9442 26753
rect 8993 26687 9060 26688
rect 9142 26193 9442 26688
rect 200 25893 9442 26193
rect 9800 31013 10100 34187
rect 10264 32192 10330 32193
rect 10264 32128 10265 32192
rect 10329 32190 10330 32192
rect 11204 32192 11270 32193
rect 11204 32190 11205 32192
rect 10329 32130 11205 32190
rect 10329 32128 10330 32130
rect 10264 32127 10330 32128
rect 11204 32128 11205 32130
rect 11269 32128 11270 32192
rect 11204 32127 11270 32128
rect 11187 31013 11253 31014
rect 9800 30949 11188 31013
rect 11252 30949 11253 31013
rect 200 20468 500 25893
rect 9552 25666 9618 25667
rect 9552 25602 9553 25666
rect 9617 25664 9618 25666
rect 9800 25664 10100 30949
rect 11187 30948 11253 30949
rect 9617 25604 10100 25664
rect 9617 25602 9618 25604
rect 9552 25601 9618 25602
rect 1280 20468 1359 20469
rect 200 20391 1281 20468
rect 1358 20391 1359 20468
rect 200 18244 500 20391
rect 1280 20390 1359 20391
rect 1292 18246 1358 18247
rect 1292 18244 1293 18246
rect 200 18184 1293 18244
rect 200 16795 500 18184
rect 1292 18182 1293 18184
rect 1357 18182 1358 18246
rect 1292 18181 1358 18182
rect 4558 16795 4727 21158
rect 9513 21003 9608 21004
rect 9800 21003 10100 25604
rect 9513 20910 9514 21003
rect 9607 20910 10100 21003
rect 9513 20909 9608 20910
rect 9800 20195 10100 20910
rect 6924 20057 10100 20195
rect 7860 19974 7920 20057
rect 8839 19982 8899 20057
rect 8836 19981 8902 19982
rect 7857 19973 7923 19974
rect 7857 19909 7858 19973
rect 7922 19909 7923 19973
rect 8836 19917 8837 19981
rect 8901 19917 8902 19981
rect 8836 19916 8902 19917
rect 7857 19908 7923 19909
rect 9800 19061 10100 20057
rect 10637 19063 10703 19064
rect 10637 19061 10638 19063
rect 9800 19001 10638 19061
rect 9800 18408 10100 19001
rect 10637 18999 10638 19001
rect 10702 18999 10703 19063
rect 10637 18998 10703 18999
rect 10370 18722 10436 18723
rect 10370 18658 10371 18722
rect 10435 18658 10436 18722
rect 10370 18657 10436 18658
rect 6850 18108 10100 18408
rect 10373 18422 10433 18657
rect 10373 18216 10689 18422
rect 200 16626 5615 16795
rect 200 16016 500 16626
rect 5446 16235 5615 16626
rect 5446 16197 9425 16235
rect 5446 16190 8307 16197
rect 5446 16126 7128 16190
rect 7192 16133 8307 16190
rect 8371 16133 9425 16197
rect 7192 16126 9425 16133
rect 5446 16066 9425 16126
rect 1340 16018 1406 16019
rect 1340 16016 1341 16018
rect 200 15956 1341 16016
rect 200 13561 500 15956
rect 1340 15954 1341 15956
rect 1405 15954 1406 16018
rect 1340 15953 1406 15954
rect 9364 15435 9430 15436
rect 9364 15371 9365 15435
rect 9429 15434 9430 15435
rect 9800 15434 10100 18108
rect 9429 15372 10100 15434
rect 9429 15371 9430 15372
rect 9364 15370 9430 15371
rect 9120 14397 9420 14398
rect 9120 14099 9121 14397
rect 9419 14099 9420 14397
rect 870 13563 936 13564
rect 870 13561 871 13563
rect 200 13501 871 13561
rect 200 2065 500 13501
rect 870 13499 871 13501
rect 935 13499 936 13563
rect 870 13498 936 13499
rect 9120 7759 9420 14099
rect 9800 13118 10100 15372
rect 10389 14399 10689 18216
rect 10388 14398 10690 14399
rect 10388 14098 10389 14398
rect 10689 14098 10690 14398
rect 10388 14097 10690 14098
rect 10533 13904 10594 14097
rect 10530 13903 10596 13904
rect 10530 13839 10531 13903
rect 10595 13839 10596 13903
rect 10530 13838 10596 13839
rect 10479 13120 10545 13121
rect 10479 13118 10480 13120
rect 9800 13058 10480 13118
rect 9604 7759 9671 7760
rect 9120 7694 9605 7759
rect 9670 7694 9671 7759
rect 9120 2065 9420 7694
rect 9604 7693 9671 7694
rect 200 1765 9420 2065
rect 9800 7216 10100 13058
rect 10479 13056 10480 13058
rect 10544 13056 10545 13120
rect 10479 13055 10545 13056
rect 10507 7217 10573 7218
rect 10507 7216 10508 7217
rect 9800 7155 10508 7216
rect 200 1000 500 1765
rect 9331 1419 9391 1765
rect 9328 1418 9394 1419
rect 9328 1354 9329 1418
rect 9393 1354 9394 1418
rect 9328 1353 9394 1354
rect 9800 894 10100 7155
rect 10507 7153 10508 7155
rect 10572 7153 10573 7217
rect 10507 7152 10573 7153
rect 11375 1635 11435 42377
rect 11572 8380 11632 43222
rect 11737 43074 11803 43075
rect 11737 43010 11738 43074
rect 11802 43010 11803 43074
rect 11737 43009 11803 43010
rect 11740 14310 11800 43009
rect 11927 20214 11987 43411
rect 21446 43279 21506 43480
rect 12087 43219 21506 43279
rect 21620 43291 21686 43292
rect 21620 43227 21621 43291
rect 21685 43227 21686 43291
rect 21620 43226 21686 43227
rect 12087 26567 12147 43219
rect 21623 43071 21683 43226
rect 12251 43011 21683 43071
rect 21801 43061 21867 43062
rect 12251 32510 12311 43011
rect 21801 42997 21802 43061
rect 21866 42997 21867 43061
rect 21801 42996 21867 42997
rect 21804 42878 21864 42996
rect 12411 42818 21864 42878
rect 12411 42753 12543 42818
rect 12411 42752 12474 42753
rect 12414 38283 12474 42752
rect 12411 38282 12477 38283
rect 12411 38218 12412 38282
rect 12476 38218 12477 38282
rect 12411 38217 12477 38218
rect 12248 32509 12314 32510
rect 12248 32445 12249 32509
rect 12313 32445 12314 32509
rect 12248 32444 12314 32445
rect 12070 26536 12162 26567
rect 12070 26472 12085 26536
rect 12149 26472 12162 26536
rect 12070 26463 12162 26472
rect 11924 20213 11990 20214
rect 11924 20149 11925 20213
rect 11989 20149 11990 20213
rect 11924 20148 11990 20149
rect 11737 14309 11803 14310
rect 11737 14245 11738 14309
rect 11802 14245 11803 14309
rect 11737 14244 11803 14245
rect 11569 8379 11635 8380
rect 11569 8315 11570 8379
rect 11634 8315 11635 8379
rect 11569 8314 11635 8315
rect 11372 1634 11438 1635
rect 11372 1570 11373 1634
rect 11437 1570 11438 1634
rect 11372 1569 11438 1570
rect 15650 894 15950 42546
rect 21946 1559 22293 43853
rect 22404 43755 22470 43756
rect 22404 43691 22405 43755
rect 22469 43753 22470 43755
rect 26558 43753 26618 45152
rect 22469 43693 26618 43753
rect 22469 43691 22470 43693
rect 22404 43690 22470 43691
rect 22391 43545 22457 43546
rect 22391 43481 22392 43545
rect 22456 43543 22457 43545
rect 27294 43543 27354 45152
rect 22456 43483 27354 43543
rect 22456 43481 22457 43483
rect 22391 43480 22457 43481
rect 22386 43291 22452 43292
rect 22386 43227 22387 43291
rect 22451 43289 22452 43291
rect 28030 43289 28090 45152
rect 22451 43229 28090 43289
rect 22451 43227 22452 43229
rect 22386 43226 22452 43227
rect 22392 43061 22458 43062
rect 22392 42997 22393 43061
rect 22457 43059 22458 43061
rect 28766 43059 28826 45152
rect 29502 44952 29562 45152
rect 30238 45087 30298 45152
rect 30173 44952 30298 45087
rect 30974 44999 31034 45152
rect 30973 44952 31034 44999
rect 31710 44952 31770 45152
rect 30173 43059 30297 44952
rect 30973 44405 31033 44952
rect 30970 44404 31036 44405
rect 30970 44340 30971 44404
rect 31035 44340 31036 44404
rect 30970 44339 31036 44340
rect 22457 42999 28826 43059
rect 22457 42997 22458 42999
rect 22392 42996 22458 42997
rect 30187 42901 30284 43059
rect 22403 42900 30284 42901
rect 22403 42805 22404 42900
rect 22499 42805 30284 42900
rect 22403 42804 30284 42805
rect 28857 894 29157 42560
rect 9800 862 29157 894
rect 9800 798 10929 862
rect 10993 798 29157 862
rect 9800 594 29157 798
rect 31282 829 31462 830
rect 31282 651 31283 829
rect 31461 651 31462 829
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 651
use psu_sequencer  psu_sequencer_0 ~/projects/adia/adia_psu_full_test/mag
timestamp 1717221846
transform 1 0 550 0 1 32800
box 0 0 9204 11348
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_0
timestamp 1717221846
transform -1 0 7798 0 1 18180
box -1786 -1640 1786 1640
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_0
timestamp 1717221846
transform 1 0 22398 0 1 3840
box -9798 -2840 9798 2840
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_1
timestamp 1717221846
transform 1 0 22398 0 1 39840
box -9798 -2840 9798 2840
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_2
timestamp 1717221846
transform 1 0 22398 0 1 33840
box -9798 -2840 9798 2840
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_3
timestamp 1717221846
transform 1 0 22398 0 1 27840
box -9798 -2840 9798 2840
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_4
timestamp 1717221846
transform 1 0 22398 0 1 21840
box -9798 -2840 9798 2840
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_5
timestamp 1717221846
transform 1 0 22398 0 1 15840
box -9798 -2840 9798 2840
use sky130_fd_pr__cap_mim_m3_1_MJ7HL7  sky130_fd_pr__cap_mim_m3_1_MJ7HL7_6
timestamp 1717221846
transform 1 0 22398 0 1 9840
box -9798 -2840 9798 2840
use sky130_fd_pr__nfet_01v8_EDB9KC  sky130_fd_pr__nfet_01v8_EDB9KC_0
timestamp 1717221846
transform 0 1 7208 -1 0 20439
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_EDB9KC  sky130_fd_pr__nfet_01v8_EDB9KC_1
timestamp 1717221846
transform 0 1 9208 -1 0 20435
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_EDB9KC  sky130_fd_pr__nfet_01v8_EDB9KC_2
timestamp 1717221846
transform 0 1 8216 -1 0 20437
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_1
timestamp 1717221846
transform -1 0 11947 0 1 13074
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_2
timestamp 1717221846
transform -1 0 11921 0 1 7175
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_3
timestamp 1717221846
transform -1 0 12047 0 1 19027
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_4
timestamp 1717221846
transform -1 0 11988 0 1 31165
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_5
timestamp 1717221846
transform -1 0 11955 0 1 25199
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_6
timestamp 1717221846
transform -1 0 12229 0 1 37059
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_8
timestamp 1717221846
transform -1 0 12127 0 1 832
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_9
timestamp 1717221846
transform -1 0 4177 0 1 19878
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_10
timestamp 1717221846
transform -1 0 4207 0 1 17664
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_EDB9KC  sky130_fd_pr__nfet_01v8_lvt_EDB9KC_11
timestamp 1717221846
transform -1 0 4197 0 1 15438
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_1
timestamp 1717221846
transform -1 0 11945 0 1 13759
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_2
timestamp 1717221846
transform -1 0 12125 0 1 1517
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_3
timestamp 1717221846
transform -1 0 12045 0 1 19712
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_4
timestamp 1717221846
transform -1 0 11986 0 1 31850
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_5
timestamp 1717221846
transform -1 0 11953 0 1 25884
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_6
timestamp 1717221846
transform -1 0 12227 0 1 37744
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_8
timestamp 1717221846
transform -1 0 11919 0 1 7860
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_9
timestamp 1717221846
transform -1 0 4175 0 1 20563
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_10
timestamp 1717221846
transform -1 0 4205 0 1 18349
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4LRBJ4  sky130_fd_pr__pfet_01v8_lvt_4LRBJ4_11
timestamp 1717221846
transform -1 0 4195 0 1 16123
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_UAQRRG  sky130_fd_pr__pfet_01v8_UAQRRG_0
timestamp 1717221846
transform 0 1 6036 -1 0 15771
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_UAQRRG  sky130_fd_pr__pfet_01v8_UAQRRG_1
timestamp 1717221846
transform 0 1 8945 -1 0 15760
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_UAQRRG  sky130_fd_pr__pfet_01v8_UAQRRG_2
timestamp 1717221846
transform 0 1 7546 -1 0 15760
box -211 -319 211 319
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717221846
transform 1 0 11394 0 1 7181
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1717221846
transform 1 0 11420 0 1 13080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1717221846
transform 1 0 5408 0 1 15304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1717221846
transform 1 0 11520 0 1 19033
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1717221846
transform 1 0 11461 0 1 31171
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1717221846
transform 1 0 11428 0 1 25205
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_7
timestamp 1717221846
transform 1 0 11702 0 1 37065
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_8
timestamp 1717221846
transform 1 0 8317 0 1 15293
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_9
timestamp 1717221846
transform 1 0 11600 0 1 838
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_10
timestamp 1717221846
transform 1 0 3650 0 1 19884
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_11
timestamp 1717221846
transform 1 0 3680 0 1 17670
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_12
timestamp 1717221846
transform 1 0 3670 0 1 15444
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_13
timestamp 1717221846
transform 1 0 6918 0 1 15293
box -38 -48 314 592
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
